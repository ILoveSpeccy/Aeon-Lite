
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f8",
X"e0738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80fb",
X"b80c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f3",
X"8f2d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f1a3",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"96e80480",
X"3d0d80fc",
X"fc087008",
X"810683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d80fc",
X"fc087008",
X"70fe0676",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80fcfc08",
X"70087081",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80fcfc08",
X"700870fd",
X"06761007",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"fcfc0870",
X"0870822c",
X"bf0683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"fcfc0870",
X"0870fe83",
X"0676822b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80fcfc08",
X"70087088",
X"2c870683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80fcfc08",
X"700870f1",
X"ff067688",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d80fcfc",
X"08700870",
X"8b2cbf06",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80fcfc",
X"08700870",
X"f88fff06",
X"768b2b07",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"fd8c0870",
X"0870882c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fd8c0870",
X"0870892c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fd8c0870",
X"08708a2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fd8c0870",
X"08708b2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"fd3d0d75",
X"81e62987",
X"2a80fcec",
X"0854730c",
X"853d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fc",
X"ce3f7280",
X"2e8338d2",
X"3f8151fc",
X"f03f8051",
X"fceb3f80",
X"51fcb83f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"9e39ff9f",
X"12519971",
X"279538d0",
X"12e01370",
X"54545189",
X"71278838",
X"8f732783",
X"38805273",
X"802e8538",
X"81801252",
X"7181ff06",
X"83e0800c",
X"853d0d04",
X"803d0d86",
X"b8c05180",
X"71708105",
X"53347086",
X"c0c02e09",
X"8106f038",
X"823d0d04",
X"fe3d0d02",
X"97053351",
X"ff863f83",
X"e0800881",
X"ff0683e0",
X"9c085452",
X"8073249b",
X"3883e0b8",
X"08137283",
X"e0bc0807",
X"53537173",
X"3483e09c",
X"08810583",
X"e09c0c84",
X"3d0d04fa",
X"3d0d8280",
X"0a1b5580",
X"57883dfc",
X"05547953",
X"74527851",
X"b5943f88",
X"3d0d04fe",
X"3d0d83e0",
X"b0085274",
X"51bbf63f",
X"83e08008",
X"8c387653",
X"755283e0",
X"b00851c7",
X"3f843d0d",
X"04fe3d0d",
X"83e0b008",
X"53755274",
X"51b6b63f",
X"83e08008",
X"8d387753",
X"765283e0",
X"b00851ff",
X"a23f843d",
X"0d04fe3d",
X"0d83e0b4",
X"0851b5aa",
X"3f83e080",
X"08818080",
X"2e098106",
X"8738b180",
X"80539a39",
X"83e0b408",
X"51b58f3f",
X"83e08008",
X"80d0802e",
X"09810692",
X"38b1b080",
X"5383e080",
X"085283e0",
X"b40851fe",
X"da3f843d",
X"0d04803d",
X"0dface3f",
X"83e08008",
X"842980fb",
X"c0057008",
X"83e0800c",
X"51823d0d",
X"04ee3d0d",
X"80438042",
X"80418070",
X"5a5bfdd4",
X"3f800b83",
X"e09c0c80",
X"0b83e0bc",
X"0c0b0b80",
X"f9fc51af",
X"fa3f8180",
X"0b83e0bc",
X"0c0b0b80",
X"fa8051af",
X"ea3f80d0",
X"0b83e09c",
X"0c783070",
X"7a078025",
X"70872b83",
X"e0bc0c51",
X"55f9b93f",
X"83e08008",
X"520b0b80",
X"fa8851af",
X"c23f80f8",
X"0b83e09c",
X"0c788132",
X"70307072",
X"07802570",
X"872b83e0",
X"bc0c5156",
X"56feeb3f",
X"83e08008",
X"520b0b80",
X"fa9451af",
X"963f81a0",
X"0b83e09c",
X"0c788232",
X"70307072",
X"07802570",
X"872b83e0",
X"bc0c5156",
X"83e0b408",
X"5256b0b1",
X"3f83e080",
X"08520b0b",
X"80fa9c51",
X"aee53f81",
X"f00b83e0",
X"9c0c810b",
X"83e0a05b",
X"5883e09c",
X"0882197a",
X"32703070",
X"72078025",
X"70872b83",
X"e0bc0c51",
X"578e3d70",
X"55ff1b54",
X"575757a4",
X"c33f7970",
X"84055b08",
X"51afe63f",
X"745483e0",
X"80085377",
X"520b0b80",
X"faa451ae",
X"963fa817",
X"83e09c0c",
X"81185877",
X"852e0981",
X"06ffae38",
X"83900b83",
X"e09c0c78",
X"87327030",
X"70720780",
X"2570872b",
X"83e0bc0c",
X"51560b0b",
X"80fab452",
X"56ade03f",
X"83e00b83",
X"e09c0c78",
X"88327030",
X"70720780",
X"2570872b",
X"83e0bc0c",
X"51560b0b",
X"80fac852",
X"56adbc3f",
X"868da051",
X"f9923f80",
X"52913d70",
X"52558ba5",
X"3f835274",
X"518b9e3f",
X"61195978",
X"80258538",
X"80599039",
X"88792585",
X"38885987",
X"39788826",
X"82ae3878",
X"822b5580",
X"f8f01508",
X"04f6e53f",
X"83e08008",
X"61575575",
X"812e0981",
X"06893883",
X"e0800810",
X"55903975",
X"ff2e0981",
X"06883883",
X"e0800881",
X"2c559075",
X"25853890",
X"55883974",
X"80248338",
X"81557451",
X"f6c23f81",
X"e339f6d5",
X"3f83e080",
X"08610555",
X"74802585",
X"38805588",
X"39877525",
X"83388755",
X"7451f6d1",
X"3f81c139",
X"60873862",
X"802e81b8",
X"38a0970b",
X"83e0d00c",
X"83e0b408",
X"518ca93f",
X"fb803f81",
X"a3396056",
X"80762598",
X"389fb60b",
X"83e0d00c",
X"83e09415",
X"70085255",
X"8c8a3f74",
X"08529139",
X"75802591",
X"3883e094",
X"150851ad",
X"a23f8052",
X"fd1951b8",
X"3962802e",
X"80ea3883",
X"e0941570",
X"0883e0a0",
X"08720c83",
X"e0a00cfd",
X"1a705351",
X"5596f93f",
X"83e08008",
X"56805196",
X"ef3f83e0",
X"80085274",
X"51938e3f",
X"75528051",
X"93873fb4",
X"3962802e",
X"af38a097",
X"0b83e0d0",
X"0c83e0b0",
X"08518ba0",
X"3f83e0b0",
X"0851acb1",
X"3f9c800a",
X"5380c080",
X"5283e080",
X"0851f99b",
X"3f81558c",
X"39628738",
X"7a802efa",
X"c5388055",
X"7483e080",
X"0c943d0d",
X"04fe3d0d",
X"f5c23f83",
X"e0800880",
X"2e863880",
X"5180f639",
X"f5ca3f83",
X"e0800880",
X"ea38f5f0",
X"3f83e080",
X"08802eaa",
X"388151f3",
X"c23f839b",
X"3f800b83",
X"e09c0cf9",
X"f43f83e0",
X"800853ff",
X"0b83e09c",
X"0c85ee3f",
X"72bd3872",
X"51f3a03f",
X"bb39f5a4",
X"3f83e080",
X"08802eb0",
X"388151f3",
X"8e3f82e7",
X"3f9fb60b",
X"83e0d00c",
X"83e0a008",
X"5189fd3f",
X"ff0b83e0",
X"9c0c85b9",
X"3f83e0a0",
X"08528051",
X"91bb3f81",
X"51f68f3f",
X"843d0d04",
X"83e08c08",
X"0283e08c",
X"0cfa3d0d",
X"800b83e0",
X"a00b83e0",
X"8c08fc05",
X"0c83e08c",
X"08f8050c",
X"aded3f83",
X"e0800886",
X"05fc0683",
X"e08c08f4",
X"050c0283",
X"e08c08f4",
X"0508310d",
X"853d7083",
X"e08c08fc",
X"05087084",
X"0583e08c",
X"08fc050c",
X"0c51aab7",
X"3f83e08c",
X"08f80508",
X"810583e0",
X"8c08f805",
X"0c83e08c",
X"08f80508",
X"862e0981",
X"06ffad38",
X"84a88080",
X"5181aa3f",
X"ff0b83e0",
X"9c0c800b",
X"83e0bc0c",
X"86b8c00b",
X"83e0b80c",
X"8151f1cb",
X"3f8151f1",
X"f43f8051",
X"f1ef3f81",
X"51f2993f",
X"8151f2f6",
X"3f8251f2",
X"c03f8e84",
X"528051a7",
X"fb3f8480",
X"805284a4",
X"808051ad",
X"d63f83e0",
X"800880d3",
X"3893d23f",
X"80fec451",
X"b2953f83",
X"e0800883",
X"e0b40854",
X"0b0b80fa",
X"d05383e0",
X"80085283",
X"e08c08f4",
X"050cace9",
X"3f83e080",
X"088438f6",
X"c13fb080",
X"805480c0",
X"80530b0b",
X"80fadc52",
X"83e08c08",
X"f4050851",
X"f6833f81",
X"51f3f33f",
X"9daa3f81",
X"51f3eb3f",
X"fccf3ffc",
X"397183e0",
X"c40c8880",
X"800b83e0",
X"c00c8480",
X"800b83e0",
X"c80c04f0",
X"3d0d80fb",
X"f4085473",
X"3383e0cc",
X"3483a080",
X"5683e0c4",
X"081683e0",
X"c0081756",
X"54743374",
X"3483e0c8",
X"08165480",
X"74348116",
X"567583a0",
X"a02e0981",
X"06db3883",
X"a4805683",
X"e0c40816",
X"83e0c008",
X"17565474",
X"33743483",
X"e0c80816",
X"54807434",
X"81165675",
X"83a4a02e",
X"098106db",
X"3883a880",
X"5683e0c4",
X"081683e0",
X"c0081756",
X"54743374",
X"3483e0c8",
X"08165480",
X"74348116",
X"567583a8",
X"902e0981",
X"06db3880",
X"fbf40854",
X"ff743480",
X"5683e0c4",
X"081683e0",
X"c8081755",
X"55733375",
X"34811656",
X"7583a080",
X"2e098106",
X"e43883b0",
X"805683e0",
X"c4081683",
X"e0c80817",
X"55557333",
X"75348116",
X"56758480",
X"802e0981",
X"06e438f2",
X"ef3f893d",
X"58a25380",
X"f9945277",
X"5180dcbc",
X"3f80578c",
X"805683e0",
X"c8081677",
X"19555573",
X"33753481",
X"16811858",
X"5676a22e",
X"098106e6",
X"3880fc98",
X"08548674",
X"3480fc9c",
X"08548074",
X"3480fc94",
X"08548074",
X"3480fc84",
X"0854af74",
X"3480fc90",
X"0854bf74",
X"3480fc8c",
X"08548074",
X"3480fc88",
X"08549f74",
X"3480fc80",
X"08548074",
X"3480fbec",
X"0854e074",
X"3480fbe4",
X"08547674",
X"3480fbe0",
X"08548374",
X"3480fbe8",
X"08548274",
X"34923d0d",
X"04fe3d0d",
X"805383e0",
X"c8081383",
X"e0c40814",
X"52527033",
X"72348113",
X"537283a0",
X"802e0981",
X"06e43883",
X"b0805383",
X"e0c80813",
X"83e0c408",
X"14525270",
X"33723481",
X"13537284",
X"80802e09",
X"8106e438",
X"83a08053",
X"83e0c808",
X"1383e0c4",
X"08145252",
X"70337234",
X"81135372",
X"83a0a02e",
X"098106e4",
X"3883a480",
X"5383e0c8",
X"081383e0",
X"c4081452",
X"52703372",
X"34811353",
X"7283a4a0",
X"2e098106",
X"e43883a8",
X"805383e0",
X"c8081383",
X"e0c40814",
X"52527033",
X"72348113",
X"537283a8",
X"902e0981",
X"06e43880",
X"fbf40851",
X"83e0cc33",
X"7134843d",
X"0d04fd3d",
X"0d755480",
X"740c800b",
X"84150c80",
X"0b88150c",
X"80fbf808",
X"70337081",
X"ff067081",
X"2a813271",
X"81327181",
X"06718106",
X"31841a0c",
X"56567083",
X"2a813271",
X"822a8132",
X"71810671",
X"81063179",
X"0c525551",
X"515180fb",
X"f0087033",
X"70098106",
X"88170c51",
X"51853d0d",
X"04fe3d0d",
X"74765452",
X"7151ff9a",
X"3f72812e",
X"a2388173",
X"268d3872",
X"822eab38",
X"72832e9f",
X"38e63971",
X"08e23884",
X"1208dd38",
X"881208d8",
X"38a03988",
X"1208812e",
X"098106cc",
X"38943988",
X"1208812e",
X"8d387108",
X"89388412",
X"08802eff",
X"b738843d",
X"0d04fc3d",
X"0d767052",
X"5580c793",
X"3f83e080",
X"0815ff05",
X"5473752e",
X"8e387333",
X"5372ae2e",
X"8638ff14",
X"54ef3977",
X"52811451",
X"80c6aa3f",
X"83e08008",
X"307083e0",
X"80080780",
X"2583e080",
X"0c53863d",
X"0d04fc3d",
X"0d767052",
X"55abfe3f",
X"83e08008",
X"54815383",
X"e0800880",
X"c1387451",
X"abc13f83",
X"e0800880",
X"fafc5383",
X"e0800852",
X"53ff8f3f",
X"83e08008",
X"a13880fb",
X"80527251",
X"ff803f83",
X"e0800892",
X"3880fb84",
X"527251fe",
X"f13f83e0",
X"8008802e",
X"83388154",
X"73537283",
X"e0800c86",
X"3d0d04fd",
X"3d0d7570",
X"5254ab9d",
X"3f815383",
X"e0800897",
X"387351aa",
X"e63f80fb",
X"885283e0",
X"800851fe",
X"b93f83e0",
X"80085372",
X"83e0800c",
X"853d0d04",
X"e03d0da3",
X"3d087052",
X"5ea18e3f",
X"83e08008",
X"33943d56",
X"54739438",
X"80fed452",
X"745184d0",
X"397d5278",
X"51a4903f",
X"84db397d",
X"51a0f63f",
X"83e08008",
X"527451a0",
X"a63f83e0",
X"d0085293",
X"3d70525b",
X"a7803f83",
X"e0800859",
X"800b83e0",
X"8008555c",
X"83e08008",
X"7c2e9438",
X"811c7452",
X"5caa813f",
X"83e08008",
X"5483e080",
X"08ee3880",
X"5aff7a43",
X"7a427a41",
X"5f790970",
X"9f2c7b06",
X"5b547b7a",
X"248438ff",
X"1c5af61a",
X"7009709f",
X"2c72067b",
X"ff125a5a",
X"52555580",
X"75259538",
X"7651a9c0",
X"3f83e080",
X"0876ff18",
X"58555773",
X"8024ed38",
X"747f2e86",
X"38ebe53f",
X"745f78ff",
X"1b70585e",
X"58807a25",
X"95387751",
X"a9963f83",
X"e0800876",
X"ff185855",
X"58738024",
X"ed38800b",
X"83e09c0c",
X"800b83e0",
X"bc0c80fb",
X"8c519deb",
X"3f81800b",
X"83e0bc0c",
X"80fb9451",
X"9ddd3fa8",
X"0b83e09c",
X"0c76802e",
X"80e43883",
X"e09c0877",
X"79327030",
X"70720780",
X"2570872b",
X"83e0bc0c",
X"51567853",
X"5656a8cd",
X"3f83e080",
X"08802e88",
X"3880fb9c",
X"519da43f",
X"7651a88f",
X"3f83e080",
X"085280fa",
X"b0519d93",
X"3f7651a8",
X"973f83e0",
X"800883e0",
X"9c085557",
X"75742586",
X"38a81656",
X"f7397583",
X"e09c0c86",
X"f07624ff",
X"98388798",
X"0b83e09c",
X"0c77802e",
X"b1387751",
X"a7cd3f83",
X"e0800878",
X"5255a7ed",
X"3f80fba4",
X"5483e080",
X"088d3887",
X"39807634",
X"fda03980",
X"fba05474",
X"53735280",
X"faec519c",
X"b23f8054",
X"80fbac51",
X"9ca93f81",
X"145473a8",
X"2e098106",
X"ef38868d",
X"a051e7f4",
X"3f805290",
X"3d705254",
X"fa873f83",
X"527351fa",
X"803f6180",
X"2e819c38",
X"7c5473ff",
X"2e963878",
X"802e819d",
X"387851a6",
X"f73f83e0",
X"8008ff15",
X"5559e739",
X"78802e81",
X"88387851",
X"a6f33f83",
X"e0800880",
X"2efc9638",
X"7851a6bb",
X"3f83e080",
X"0883e080",
X"085380fa",
X"f45254bf",
X"e33f83e0",
X"8008a538",
X"7a5180c1",
X"9a3f83e0",
X"80085574",
X"ff165654",
X"807425fb",
X"fd38741b",
X"70335556",
X"73af2efe",
X"cc38e839",
X"7a5180c0",
X"f63f8253",
X"80faf852",
X"83e08008",
X"1b5180d2",
X"9b3f7a51",
X"80c0e03f",
X"735283e0",
X"80081b51",
X"80c0b83f",
X"fbc4397f",
X"88296010",
X"057a0561",
X"055afbf5",
X"39a23d0d",
X"04803d0d",
X"81ff5180",
X"0b83e0dc",
X"1234ff11",
X"5170f438",
X"823d0d04",
X"ff3d0d73",
X"70335351",
X"81113371",
X"34718112",
X"34833d0d",
X"04fb3d0d",
X"77795656",
X"80707155",
X"55527175",
X"25ac3872",
X"16703370",
X"147081ff",
X"06555151",
X"51717427",
X"89388112",
X"7081ff06",
X"53517181",
X"147083ff",
X"ff065552",
X"54747324",
X"d6387183",
X"e0800c87",
X"3d0d04fd",
X"3d0d7554",
X"948f3f83",
X"e0800880",
X"2ef63883",
X"e2f80886",
X"057081ff",
X"06525391",
X"e83f8439",
X"eef33f93",
X"f03f83e0",
X"8008812e",
X"f33892cb",
X"3f83e080",
X"08743492",
X"c23f83e0",
X"80088115",
X"3492b83f",
X"83e08008",
X"82153492",
X"ae3f83e0",
X"80088315",
X"3492a43f",
X"83e08008",
X"84153484",
X"39eeb23f",
X"93af3f83",
X"e0800880",
X"2ef33873",
X"3383e0dc",
X"34811433",
X"83e0dd34",
X"82143383",
X"e0de3483",
X"143383e0",
X"df348452",
X"83e0dc51",
X"fea73f83",
X"e0800881",
X"ff068415",
X"33555372",
X"742e0981",
X"068c3892",
X"a03f83e0",
X"8008802e",
X"9a3883e2",
X"f808a82e",
X"09810689",
X"38860b83",
X"e2f80c87",
X"39a80b83",
X"e2f80c80",
X"e451e3ec",
X"3f853d0d",
X"04f43d0d",
X"7e605955",
X"805d8075",
X"822b7183",
X"e2fc120c",
X"83e39017",
X"5b5b5776",
X"79347777",
X"2e83b138",
X"76527751",
X"9be13f8e",
X"3dfc0554",
X"905383e2",
X"e4527751",
X"9b983f7c",
X"5675902e",
X"09810683",
X"8f3883e2",
X"e451fd84",
X"3f83e2e6",
X"51fcfd3f",
X"83e2e851",
X"fcf63f76",
X"83e2f40c",
X"775198e5",
X"3f80fb80",
X"5283e080",
X"0851f5ea",
X"3f83e080",
X"08812e09",
X"810680d3",
X"387683e3",
X"8c0c820b",
X"83e2e434",
X"ff960b83",
X"e2e53477",
X"519bab3f",
X"83e08008",
X"5583e080",
X"08772588",
X"3883e080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"e2e63474",
X"83e2e734",
X"7683e2e8",
X"34ff800b",
X"83e2e934",
X"818f3983",
X"e2e43383",
X"e2e53371",
X"882b0756",
X"5b7483ff",
X"ff2e0981",
X"0680e738",
X"fe800b83",
X"e38c0c81",
X"0b83e2f4",
X"0cff0b83",
X"e2e434ff",
X"0b83e2e5",
X"3477519a",
X"b93f83e0",
X"800883e3",
X"940c83e0",
X"80085583",
X"e0800880",
X"25883883",
X"e080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583e2e6",
X"347483e2",
X"e7347683",
X"e2e834ff",
X"800b83e2",
X"e934810b",
X"83e2f334",
X"a4397485",
X"962e0981",
X"0680fd38",
X"7583e38c",
X"0c775199",
X"ee3f83e2",
X"f33383e0",
X"80080755",
X"7483e2f3",
X"3483e2f3",
X"33810655",
X"74802e83",
X"38845783",
X"e2e83383",
X"e2e93371",
X"882b0756",
X"5c748180",
X"2e098106",
X"a13883e2",
X"e63383e2",
X"e7337188",
X"2b07565b",
X"ad807527",
X"87387682",
X"07579c39",
X"76810757",
X"96397482",
X"802e0981",
X"06873876",
X"83075787",
X"397481ff",
X"268a3877",
X"83e2fc1b",
X"0c767934",
X"8e3d0d04",
X"803d0d72",
X"842983e2",
X"fc057008",
X"83e0800c",
X"51823d0d",
X"04fe3d0d",
X"800b83e2",
X"e00c800b",
X"83e2dc0c",
X"ff0b83e0",
X"d80ca80b",
X"83e2f80c",
X"ae518ca5",
X"3f800b83",
X"e2fc5452",
X"80737084",
X"05550c81",
X"12527184",
X"2e098106",
X"ef38843d",
X"0d04fe3d",
X"0d740284",
X"05960522",
X"53537180",
X"2e963872",
X"70810554",
X"33518cc4",
X"3fff1270",
X"83ffff06",
X"5152e739",
X"843d0d04",
X"fe3d0d02",
X"92052253",
X"82ac51df",
X"873f80c3",
X"518ca13f",
X"819651de",
X"fb3f7252",
X"83e0dc51",
X"ffb43f72",
X"5283e0dc",
X"51f8e63f",
X"83e08008",
X"81ff0651",
X"8bfe3f84",
X"3d0d04ff",
X"b13d0d80",
X"d13df805",
X"51f9903f",
X"83e2e008",
X"810583e2",
X"e00c80cf",
X"3d33cf11",
X"7081ff06",
X"51565674",
X"832688cd",
X"38758f06",
X"ff055675",
X"83e0d808",
X"2e9b3875",
X"83269638",
X"7583e0d8",
X"0c758429",
X"83e2fc05",
X"70085355",
X"7551faa1",
X"3f807624",
X"88a93875",
X"842983e2",
X"fc055574",
X"08802e88",
X"9a3883e0",
X"d8088429",
X"83e2fc05",
X"70080288",
X"0582b905",
X"33525b55",
X"7480d22e",
X"849a3874",
X"80d22490",
X"3874bf2e",
X"9c387480",
X"d02e81d1",
X"3887d939",
X"7480d32e",
X"80cf3874",
X"80d72e81",
X"c03887c8",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055656",
X"8b803f80",
X"c1518ab4",
X"3ff6e23f",
X"860b83e0",
X"dc348152",
X"83e0dc51",
X"8bef3f81",
X"51fde93f",
X"74893886",
X"0b83e2f8",
X"0c8739a8",
X"0b83e2f8",
X"0c8acf3f",
X"80c1518a",
X"833ff6b1",
X"3f900b83",
X"e2f33381",
X"06565674",
X"802e8338",
X"985683e2",
X"e83383e2",
X"e9337188",
X"2b075659",
X"7481802e",
X"0981069c",
X"3883e2e6",
X"3383e2e7",
X"3371882b",
X"075657ad",
X"8075278c",
X"38758180",
X"07568539",
X"75a00756",
X"7583e0dc",
X"34ff0b83",
X"e0dd34e0",
X"0b83e0de",
X"34800b83",
X"e0df3484",
X"5283e0dc",
X"518ae63f",
X"84518686",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055659",
X"89c43f79",
X"5194c03f",
X"83e08008",
X"802e8a38",
X"80ce5188",
X"eb3f85dd",
X"3980c151",
X"88e23f89",
X"ea3f87ee",
X"3f83e38c",
X"08588375",
X"259b3883",
X"e2e83383",
X"e2e93371",
X"882b07fc",
X"1771297a",
X"05838005",
X"5a51578d",
X"39748180",
X"2918ff80",
X"05588180",
X"57805676",
X"762e9238",
X"88c13f83",
X"e0800883",
X"e0dc1734",
X"811656eb",
X"3988b03f",
X"83e08008",
X"81ff0677",
X"5383e0dc",
X"5256f4dd",
X"3f83e080",
X"0881ff06",
X"5575752e",
X"09810681",
X"843888b2",
X"3f80c151",
X"87e63f88",
X"ee3f7752",
X"795192df",
X"3f805e80",
X"d13dfdf4",
X"05547653",
X"83e0dc52",
X"795190e8",
X"3f0282b9",
X"05335581",
X"587480d7",
X"2e098106",
X"bc3880d1",
X"3dfdf005",
X"5476538f",
X"3d70537a",
X"525991ee",
X"3f805676",
X"762ea238",
X"751983e0",
X"dc173371",
X"33707232",
X"70307080",
X"2570307e",
X"06811d5d",
X"5e515151",
X"525b55db",
X"3982ac51",
X"d9d63f77",
X"802e8638",
X"80c35184",
X"3980ce51",
X"86e63f87",
X"ee3f85f2",
X"3f83d539",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"05595580",
X"705d5987",
X"893f80c1",
X"5186bd3f",
X"83e2f408",
X"792e82db",
X"3883e394",
X"0880fc05",
X"5580fd52",
X"7451bdc1",
X"3f83e080",
X"085b7782",
X"24b238ff",
X"1870872b",
X"83ffff80",
X"0680fd90",
X"0583e0dc",
X"59575581",
X"80557570",
X"81055733",
X"77708105",
X"5934ff15",
X"7081ff06",
X"515574ea",
X"38828a39",
X"7782e82e",
X"81aa3877",
X"82e92e09",
X"810681b1",
X"3880fba8",
X"518cd43f",
X"78587787",
X"32703070",
X"72078025",
X"7a8a3270",
X"30707207",
X"80257307",
X"53545a51",
X"57557580",
X"2e973878",
X"78269238",
X"a00b83e0",
X"dc1a3481",
X"197081ff",
X"065a55eb",
X"39811870",
X"81ff0659",
X"558a7827",
X"ffbc388f",
X"5883e0d7",
X"183383e0",
X"dc1934ff",
X"187081ff",
X"06595577",
X"8426ea38",
X"9058800b",
X"83e0dc19",
X"34811870",
X"81ff0670",
X"982b5259",
X"55748025",
X"e93880c6",
X"557a858f",
X"24843880",
X"c2557483",
X"e0dc3480",
X"f10b83e0",
X"df34810b",
X"83e0e034",
X"7a83e0dd",
X"347a882c",
X"557483e0",
X"de3480c9",
X"3982f078",
X"2580c238",
X"7780fd29",
X"fd97d305",
X"5279518f",
X"963f80d1",
X"3dfdec05",
X"5480fd53",
X"83e0dc52",
X"79518eca",
X"3f7b8119",
X"59567580",
X"fc248338",
X"78587788",
X"2c557483",
X"e1d93477",
X"83e1da34",
X"7583e1db",
X"34818059",
X"80ca3983",
X"e38c0857",
X"8378259b",
X"3883e2e8",
X"3383e2e9",
X"3371882b",
X"07fc1a71",
X"29790583",
X"80055951",
X"598d3977",
X"81802917",
X"ff800557",
X"81805976",
X"5279518e",
X"a63f80d1",
X"3dfdec05",
X"54785383",
X"e0dc5279",
X"518ddb3f",
X"7851f6d8",
X"3f84943f",
X"82983f8b",
X"3983e2dc",
X"08810583",
X"e2dc0c80",
X"d13d0d04",
X"f6f93fdf",
X"a83ff939",
X"fc3d0d76",
X"78718429",
X"83e2fc05",
X"70085153",
X"5353709e",
X"3880ce72",
X"3480cf0b",
X"81133480",
X"ce0b8213",
X"3480c50b",
X"83133470",
X"84133480",
X"e73983e3",
X"90133354",
X"80d27234",
X"73822a70",
X"81065151",
X"80cf5370",
X"843880d7",
X"53728113",
X"34a00b82",
X"13347383",
X"06517081",
X"2e9e3870",
X"81248838",
X"70802e8f",
X"389f3970",
X"822e9238",
X"70832e92",
X"38933980",
X"d8558e39",
X"80d35589",
X"3980cd55",
X"843980c4",
X"55748313",
X"3480c40b",
X"84133480",
X"0b851334",
X"863d0d04",
X"fe3d0d80",
X"fca80870",
X"337081ff",
X"0670842a",
X"81328106",
X"55515253",
X"71802e8c",
X"38a87334",
X"80fca808",
X"51b87134",
X"7183e080",
X"0c843d0d",
X"04fe3d0d",
X"80fca808",
X"70337081",
X"ff067085",
X"2a813281",
X"06555152",
X"5371802e",
X"8c389873",
X"3480fca8",
X"0851b871",
X"347183e0",
X"800c843d",
X"0d04803d",
X"0d80fca4",
X"08519371",
X"3480fcb0",
X"0851ff71",
X"34823d0d",
X"04fe3d0d",
X"02930533",
X"80fca408",
X"53538072",
X"348a51d3",
X"a33fd33f",
X"80fcb408",
X"5280f872",
X"3480fccc",
X"08528072",
X"34fa1380",
X"fcd40853",
X"53727234",
X"80fcbc08",
X"52807234",
X"80fcc408",
X"52727234",
X"80fca808",
X"52807234",
X"80fca808",
X"52b87234",
X"843d0d04",
X"ff3d0d02",
X"8f053380",
X"fcac0852",
X"52717134",
X"fe9e3f83",
X"e0800880",
X"2ef63883",
X"3d0d0480",
X"3d0d8439",
X"dc933ffe",
X"b83f83e0",
X"8008802e",
X"f33880fc",
X"ac087033",
X"7081ff06",
X"83e0800c",
X"5151823d",
X"0d04803d",
X"0d80fca4",
X"0851a371",
X"3480fcb0",
X"0851ff71",
X"3480fca8",
X"0851a871",
X"3480fca8",
X"0851b871",
X"34823d0d",
X"04803d0d",
X"80fca408",
X"70337081",
X"c0067030",
X"70802583",
X"e0800c51",
X"51515182",
X"3d0d04ff",
X"3d0d80fc",
X"a8087033",
X"7081ff06",
X"70832a81",
X"32708106",
X"51515152",
X"5270802e",
X"e538b072",
X"3480fca8",
X"0851b871",
X"34833d0d",
X"04803d0d",
X"80fce008",
X"70088106",
X"83e0800c",
X"51823d0d",
X"04fd3d0d",
X"75775454",
X"80732594",
X"38737081",
X"05553352",
X"80fbb051",
X"859d3fff",
X"1353e939",
X"853d0d04",
X"f63d0d7c",
X"7e60625a",
X"5d5b5680",
X"59815585",
X"39747a29",
X"55745275",
X"51b5923f",
X"83e08008",
X"7a27ee38",
X"74802e80",
X"dd387452",
X"7551b4fd",
X"3f83e080",
X"08755376",
X"5254b5a4",
X"3f83e080",
X"087a5375",
X"5256b4e5",
X"3f83e080",
X"08793070",
X"7b079f2a",
X"70778024",
X"07515154",
X"55728738",
X"83e08008",
X"c5387681",
X"18b01655",
X"58588974",
X"258b38b7",
X"14537a85",
X"3880d714",
X"53727834",
X"811959ff",
X"9f398077",
X"348c3d0d",
X"04f73d0d",
X"7b7d7f62",
X"029005bb",
X"05335759",
X"565a5ab0",
X"58728338",
X"a0587570",
X"70810552",
X"33715954",
X"55903980",
X"74258e38",
X"ff147770",
X"81055933",
X"545472ef",
X"3873ff15",
X"55538073",
X"25893877",
X"52795178",
X"2def3975",
X"33755753",
X"72802e90",
X"38725279",
X"51782d75",
X"70810557",
X"3353ed39",
X"8b3d0d04",
X"ee3d0d64",
X"66696970",
X"70810552",
X"335b4a5c",
X"5e5e7680",
X"2e82f938",
X"76a52e09",
X"810682e0",
X"38807041",
X"67707081",
X"05523371",
X"4a59575f",
X"76b02e09",
X"81068c38",
X"75708105",
X"57337648",
X"57815fd0",
X"17567589",
X"2680da38",
X"76675c59",
X"805c9339",
X"778a2480",
X"c3387b8a",
X"29187b70",
X"81055d33",
X"5a5cd019",
X"7081ff06",
X"58588977",
X"27a438ff",
X"9f197081",
X"ff06ffa9",
X"1b5a5156",
X"85762792",
X"38ffbf19",
X"7081ff06",
X"51567585",
X"268a38c9",
X"19587780",
X"25ffb938",
X"7a477b40",
X"7881ff06",
X"577680e4",
X"2e80e538",
X"7680e424",
X"a7387680",
X"d82e8186",
X"387680d8",
X"24903876",
X"802e81cc",
X"3876a52e",
X"81b63881",
X"b9397680",
X"e32e818c",
X"3881af39",
X"7680f52e",
X"9b387680",
X"f5248b38",
X"7680f32e",
X"81813881",
X"99397680",
X"f82e80ca",
X"38818f39",
X"913d7055",
X"5780538a",
X"5279841b",
X"7108535b",
X"56fc813f",
X"7655ab39",
X"79841b71",
X"08943d70",
X"5b5b525b",
X"56758025",
X"8c387530",
X"56ad7834",
X"0280c105",
X"57765480",
X"538a5275",
X"51fbd53f",
X"77557e54",
X"b839913d",
X"70557780",
X"d8327030",
X"70802556",
X"51585690",
X"5279841b",
X"7108535b",
X"57fbb13f",
X"7555db39",
X"79841b83",
X"1233545b",
X"56983979",
X"841b7108",
X"575b5680",
X"547f537c",
X"527d51fc",
X"9c3f8739",
X"76527d51",
X"7c2d6670",
X"33588105",
X"47fd8339",
X"943d0d04",
X"7283e090",
X"0c7183e0",
X"940c04fb",
X"3d0d883d",
X"70708405",
X"52085754",
X"755383e0",
X"90085283",
X"e0940851",
X"fcc63f87",
X"3d0d04ff",
X"3d0d7370",
X"08535102",
X"93053372",
X"34700881",
X"05710c83",
X"3d0d04fc",
X"3d0d873d",
X"88115578",
X"5480c0c3",
X"5351fc98",
X"3f805287",
X"3d51d03f",
X"863d0d04",
X"fd3d0d75",
X"705254a5",
X"8e3f83e0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83e0",
X"8008732e",
X"a13883e0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183e0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83e5bc08",
X"248a38a5",
X"f83fff0b",
X"83e5bc0c",
X"800b83e0",
X"800c04ff",
X"3d0d7352",
X"83e39808",
X"722e8d38",
X"d93f7151",
X"97853f71",
X"83e3980c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088191",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883e5ec",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83e5bc08",
X"2e8438ff",
X"893f83e5",
X"bc088025",
X"a6387589",
X"2b5199f1",
X"3f83e5ec",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5197d63f",
X"761483e5",
X"ec0c7583",
X"e5bc0c74",
X"53765278",
X"51a4a93f",
X"83e08008",
X"83e5ec08",
X"1683e5ec",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383e0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe9b3f",
X"7651feaf",
X"3f863dfc",
X"055302a2",
X"05225277",
X"5196f63f",
X"79863d22",
X"710c5483",
X"e0800854",
X"83e08008",
X"802e8338",
X"81547383",
X"e0800c86",
X"3d0d04fd",
X"3d0d7683",
X"e5bc0853",
X"53807224",
X"89387173",
X"2e8438fd",
X"d13f7551",
X"fde53f72",
X"5198be3f",
X"73527380",
X"2e833881",
X"527183e0",
X"800c853d",
X"0d04803d",
X"0d7280c0",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d72bc",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"c40b83e0",
X"800c04fd",
X"3d0d7577",
X"71547053",
X"5553a0e7",
X"3f82c813",
X"08bc150c",
X"82c01308",
X"80c0150c",
X"fcec3f73",
X"5194983f",
X"7383e398",
X"0c83e080",
X"085383e0",
X"8008802e",
X"83388153",
X"7283e080",
X"0c853d0d",
X"04fd3d0d",
X"75775553",
X"fcc03f72",
X"802ea538",
X"bc130852",
X"73519ff1",
X"3f83e080",
X"088f3877",
X"527251ff",
X"9a3f83e0",
X"8008538a",
X"3982cc13",
X"0853d839",
X"81537283",
X"e0800c85",
X"3d0d04fe",
X"3d0dff0b",
X"83e5bc0c",
X"7483e39c",
X"0c7583e5",
X"b80ca0de",
X"3f83e080",
X"0881ff06",
X"52815371",
X"993883e5",
X"d4518f90",
X"3f83e080",
X"085283e0",
X"8008802e",
X"83387252",
X"71537283",
X"e0800c84",
X"3d0d04fa",
X"3d0d787a",
X"82c41208",
X"82c41208",
X"70722459",
X"56565757",
X"73732e09",
X"81069138",
X"80c01652",
X"80c01751",
X"9de23f83",
X"e0800855",
X"7483e080",
X"0c883d0d",
X"04f63d0d",
X"7c5b807b",
X"715c5457",
X"7a772e8c",
X"38811a82",
X"cc140854",
X"5a72f638",
X"805980d9",
X"397a5481",
X"5780707b",
X"7b315a57",
X"55ff1853",
X"74732580",
X"c13882cc",
X"14085273",
X"51ff8c3f",
X"800b83e0",
X"800825a1",
X"3882cc14",
X"0882cc11",
X"0882cc16",
X"0c7482cc",
X"120c5375",
X"802e8638",
X"7282cc17",
X"0c725480",
X"577382cc",
X"15088117",
X"575556ff",
X"b8398119",
X"59800bff",
X"1b545478",
X"73258338",
X"81547681",
X"32707506",
X"515372ff",
X"90388c3d",
X"0d04f73d",
X"0d7b7d5a",
X"5a82d052",
X"83e5b808",
X"51a89e3f",
X"83e08008",
X"57f9e33f",
X"795283e5",
X"c05196c7",
X"3f83e080",
X"08538054",
X"83e08008",
X"742e0981",
X"06828338",
X"83e39c08",
X"0b0b80fa",
X"f4537052",
X"559da03f",
X"0b0b80fa",
X"f45280c0",
X"15519d93",
X"3f74bc16",
X"0c7282c0",
X"160c810b",
X"82c4160c",
X"810b82c8",
X"160cff17",
X"73575781",
X"973983e3",
X"a8337082",
X"2a708106",
X"51545472",
X"81863873",
X"812a8106",
X"587780fc",
X"3876802e",
X"81903882",
X"d015ff18",
X"75842a81",
X"0682c413",
X"0c83e3a8",
X"33810682",
X"c8130c7b",
X"54715358",
X"569cb43f",
X"75519ccb",
X"3f83e080",
X"081653af",
X"73708105",
X"553472bc",
X"170c83e3",
X"a9527251",
X"9c953f83",
X"e3a00882",
X"c0170c83",
X"e3b65283",
X"9015519c",
X"823f7782",
X"cc170c78",
X"802e8d38",
X"7551782d",
X"83e08008",
X"802e8d38",
X"74802e86",
X"387582cc",
X"160c7555",
X"83e3a052",
X"83e5c051",
X"95e73f83",
X"e080088a",
X"3883e3a9",
X"335372fe",
X"d138800b",
X"82cc170c",
X"78802e89",
X"3883e39c",
X"0851fcb9",
X"3f83e39c",
X"08547383",
X"e0800c8b",
X"3d0d04ff",
X"3d0d8052",
X"7351fdb6",
X"3f833d0d",
X"04f03d0d",
X"62705254",
X"f6923f83",
X"e0800874",
X"53873d70",
X"535555f6",
X"b23ff792",
X"3f7351d3",
X"3f635374",
X"5283e080",
X"0851fab9",
X"3f923d0d",
X"047183e0",
X"800c0480",
X"c01283e0",
X"800c0480",
X"3d0d7282",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"82cc1108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"7282c411",
X"0883e080",
X"0c51823d",
X"0d04f63d",
X"0d7c83e0",
X"98085959",
X"81792782",
X"a9387888",
X"19082782",
X"a1387733",
X"5675822e",
X"819b3875",
X"82248938",
X"75812e8d",
X"38828b39",
X"75832e81",
X"b7388282",
X"397883ff",
X"ff067081",
X"2a117083",
X"ffff0670",
X"83ff0671",
X"892a903d",
X"5f525a51",
X"51557683",
X"ff2e8e38",
X"82547653",
X"8c180815",
X"527951a9",
X"39755476",
X"538c1808",
X"15527951",
X"9ad83f83",
X"e0800881",
X"bd387554",
X"83e08008",
X"538c1808",
X"15810552",
X"8c3dfd05",
X"519abb3f",
X"83e08008",
X"81a03802",
X"a905338c",
X"3d337188",
X"2b077a81",
X"0671842a",
X"53575856",
X"74863876",
X"9fff0656",
X"75558180",
X"39755478",
X"1083fe06",
X"5378882a",
X"8c190805",
X"528c3dfc",
X"055199fa",
X"3f83e080",
X"0880df38",
X"02a90533",
X"8c3d3371",
X"882b0756",
X"5780d139",
X"84547882",
X"2b83fc06",
X"5378872a",
X"8c190805",
X"528c3dfc",
X"055199ca",
X"3f83e080",
X"08b03802",
X"ab053302",
X"8405aa05",
X"3371982b",
X"71902b07",
X"028c05a9",
X"05337088",
X"2b720790",
X"3d337180",
X"fffffe80",
X"06075152",
X"53575856",
X"83398155",
X"7483e080",
X"0c8c3d0d",
X"04fb3d0d",
X"83e09808",
X"fe198812",
X"08fe0555",
X"56548056",
X"7473278d",
X"38821433",
X"75712994",
X"16080557",
X"537583e0",
X"800c873d",
X"0d04fc3d",
X"0d7683e0",
X"98085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"ff933f83",
X"e0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183e080",
X"0c863d0d",
X"04fa3d0d",
X"7883e098",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fbdb3f",
X"81527183",
X"e0800827",
X"a8388352",
X"83e08008",
X"88170827",
X"9c3883e0",
X"80088c16",
X"0c83e080",
X"0851fdf9",
X"3f83e080",
X"0890160c",
X"73752380",
X"527183e0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585d5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"a0269138",
X"7a51fdd2",
X"3f83e080",
X"0856807c",
X"3483a839",
X"933d841c",
X"0870585a",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"38807059",
X"5d887f08",
X"5f5a7c81",
X"1e7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535f57",
X"557480d8",
X"3876ae2e",
X"09810683",
X"38815577",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675ac",
X"3888588b",
X"5affab39",
X"ff9f1755",
X"74992689",
X"38e01770",
X"81ff0658",
X"55778119",
X"7081ff06",
X"721c535a",
X"57557675",
X"34ff8739",
X"7c1e7f0c",
X"805576a0",
X"26833881",
X"55748b1a",
X"347a51fc",
X"913f83e0",
X"800880f5",
X"38a0547a",
X"2270852b",
X"83e00654",
X"55901b08",
X"527b5194",
X"d13f83e0",
X"80085783",
X"e0800881",
X"82387b33",
X"5574802e",
X"80f5388b",
X"1c337083",
X"2a708106",
X"51565674",
X"b4388b7c",
X"841d0883",
X"e0800859",
X"5b5b58ff",
X"185877ff",
X"2e9a3879",
X"7081055b",
X"33797081",
X"055b3371",
X"71315256",
X"5675802e",
X"e2388639",
X"75802ebc",
X"387a51fb",
X"f43fff86",
X"3983e080",
X"085683e0",
X"8008802e",
X"a93883e0",
X"8008832e",
X"09810680",
X"de38841b",
X"088b1133",
X"51557480",
X"d2388456",
X"80cd3983",
X"56ec3981",
X"5680c439",
X"7656841b",
X"088b1133",
X"515574b7",
X"388b1c33",
X"70842a70",
X"81065156",
X"5774802e",
X"d538951c",
X"33941d33",
X"71982b71",
X"902b079b",
X"1f337f9a",
X"05337188",
X"2b077207",
X"7f88050c",
X"5a585658",
X"fcda3975",
X"83e0800c",
X"903d0d04",
X"f83d0d7a",
X"7c595782",
X"5483fe53",
X"77527651",
X"92e03f83",
X"5683e080",
X"0880ec38",
X"81173377",
X"3371882b",
X"07565682",
X"567482d4",
X"d52e0981",
X"0680d438",
X"7554b653",
X"77527651",
X"92b43f83",
X"e0800898",
X"38811733",
X"77337188",
X"2b0783e0",
X"80085256",
X"56748182",
X"c62eac38",
X"825480d2",
X"53775276",
X"51928b3f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62e83",
X"38815675",
X"83e0800c",
X"8a3d0d04",
X"ec3d0d66",
X"59800b83",
X"e0980c78",
X"5678802e",
X"83e83891",
X"a53f83e0",
X"80088106",
X"55825674",
X"83d83874",
X"75538e3d",
X"70535858",
X"fec23f83",
X"e0800881",
X"ff065675",
X"812e0981",
X"0680d438",
X"905483be",
X"53745276",
X"5191973f",
X"83e08008",
X"80c9388e",
X"3d335574",
X"802e80c9",
X"3802bb05",
X"33028405",
X"ba053371",
X"982b7190",
X"2b07028c",
X"05b90533",
X"70882b72",
X"07943d33",
X"71077058",
X"7c575452",
X"5d575956",
X"fde63f83",
X"e0800881",
X"ff065675",
X"832e0981",
X"06863881",
X"5682db39",
X"75802e86",
X"38875682",
X"d139a454",
X"8d537752",
X"765190ae",
X"3f815683",
X"e0800882",
X"bd3802ba",
X"05330284",
X"05b90533",
X"71882b07",
X"585c76ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"0754525d",
X"57585602",
X"b3053377",
X"71290288",
X"05b20533",
X"028c05b1",
X"05337188",
X"2b07701c",
X"708c1f0c",
X"5e595758",
X"5c8d3d33",
X"821a3402",
X"b505338f",
X"3d337188",
X"2b07595b",
X"77841a23",
X"02b70533",
X"028405b6",
X"05337188",
X"2b07565b",
X"74ab3802",
X"80c60533",
X"02840580",
X"c5053371",
X"982b7190",
X"2b07953d",
X"3370882b",
X"72070294",
X"0580c305",
X"33710751",
X"5253575d",
X"5b747631",
X"77317884",
X"2a8f3d33",
X"54717131",
X"53565698",
X"803f83e0",
X"80088205",
X"70881b0c",
X"709ff626",
X"81055755",
X"83fff675",
X"27833883",
X"56757934",
X"75832e09",
X"8106af38",
X"0280d205",
X"33028405",
X"80d10533",
X"71982b71",
X"902b0798",
X"3d337088",
X"2b720702",
X"940580cf",
X"05337107",
X"901f0c52",
X"5d575956",
X"8639761a",
X"901a0c84",
X"19228c1a",
X"08187184",
X"2a05941b",
X"0c5c800b",
X"811a3478",
X"83e0980c",
X"80567583",
X"e0800c96",
X"3d0d04e9",
X"3d0d83e0",
X"98085686",
X"5475802e",
X"81a63880",
X"0b811734",
X"993de011",
X"466a54c0",
X"1153ec05",
X"51f6cf3f",
X"83e08008",
X"5483e080",
X"08818538",
X"893d3354",
X"73802e93",
X"3802ab05",
X"3370842a",
X"70810651",
X"55557380",
X"2e863883",
X"5480e539",
X"02b50533",
X"8f3d3371",
X"982b7190",
X"2b07028c",
X"05bb0533",
X"029005ba",
X"05337188",
X"2b077207",
X"a01b0c02",
X"9005bf05",
X"33029405",
X"be053371",
X"982b7190",
X"2b07029c",
X"05bd0533",
X"70882b72",
X"07993d33",
X"71077f9c",
X"050c5283",
X"e0800898",
X"1f0c565a",
X"52525357",
X"5957810b",
X"81173483",
X"e0800854",
X"7383e080",
X"0c993d0d",
X"04f53d0d",
X"7d600288",
X"05ba0522",
X"7283e098",
X"085b5d5a",
X"5c5c807b",
X"23865676",
X"802e81e0",
X"38811733",
X"81065585",
X"5674802e",
X"81d2389c",
X"17089818",
X"08315574",
X"78278738",
X"7483ffff",
X"06587780",
X"2e81ae38",
X"98170870",
X"83ff0656",
X"567480ca",
X"38821733",
X"ff057689",
X"2a067081",
X"ff065a55",
X"78a03875",
X"8738a017",
X"08558d39",
X"a4170851",
X"efe03f83",
X"e0800855",
X"81752780",
X"f83874a4",
X"180ca417",
X"0851f28d",
X"3f83e080",
X"08802e80",
X"e43883e0",
X"800819a8",
X"180c9817",
X"0883ff06",
X"84807131",
X"7083ffff",
X"06585155",
X"77762783",
X"38775675",
X"54981708",
X"83ff0653",
X"a8170852",
X"79557b83",
X"387b5574",
X"518ad33f",
X"83e08008",
X"a4389817",
X"08169818",
X"0c751a78",
X"77317083",
X"ffff067d",
X"22790552",
X"5a565a74",
X"7b23fece",
X"39805688",
X"39800b81",
X"18348156",
X"7583e080",
X"0c8d3d0d",
X"04fa3d0d",
X"7883e098",
X"08555686",
X"5573802e",
X"81dc3881",
X"14338106",
X"53855572",
X"802e81ce",
X"389c1408",
X"53727627",
X"83387256",
X"98140857",
X"800b9815",
X"0c75802e",
X"81a93882",
X"14337089",
X"2b565376",
X"802eb538",
X"7452ff16",
X"5192ee3f",
X"83e08008",
X"ff187654",
X"70535853",
X"92df3f83",
X"e0800873",
X"26963874",
X"30707806",
X"7098170c",
X"777131a4",
X"17085258",
X"51538939",
X"a0140870",
X"a4160c53",
X"747627b4",
X"387251ed",
X"c13f83e0",
X"80085381",
X"0b83e080",
X"082780cb",
X"3883e080",
X"08881508",
X"2780c038",
X"83e08008",
X"a4150c98",
X"14081598",
X"150c7575",
X"3156c939",
X"98140816",
X"7098160c",
X"735256ef",
X"c83f83e0",
X"8008802e",
X"96388214",
X"33ff0576",
X"892a0683",
X"e0800805",
X"a8150c80",
X"55883980",
X"0b811534",
X"81557483",
X"e0800c88",
X"3d0d04ee",
X"3d0d6456",
X"865583e0",
X"9808802e",
X"80f63894",
X"3df41184",
X"180c6654",
X"d4055275",
X"51f1973f",
X"83e08008",
X"5583e080",
X"0880cf38",
X"893d3354",
X"73802ebc",
X"3802ab05",
X"3370842a",
X"70810651",
X"55558455",
X"73802ebc",
X"3802b505",
X"338f3d33",
X"71982b71",
X"902b0702",
X"8c05bb05",
X"33029005",
X"ba053371",
X"882b0772",
X"07881b0c",
X"53575957",
X"7551eed2",
X"3f83e080",
X"08557483",
X"2e098106",
X"83388455",
X"7483e080",
X"0c943d0d",
X"04e43d0d",
X"6ea13d08",
X"405d8656",
X"83e09808",
X"802e849b",
X"389e3df4",
X"05841e0c",
X"7e98387c",
X"51ee973f",
X"83e08008",
X"56848439",
X"81418280",
X"39834181",
X"fb39933d",
X"7f960541",
X"59807f82",
X"95055f56",
X"756081ff",
X"05348341",
X"901d0876",
X"2e81dd38",
X"a0547c22",
X"70852b83",
X"e0065458",
X"901d0852",
X"785186ae",
X"3f83e080",
X"084183e0",
X"8008ffb8",
X"3878335c",
X"7b802eff",
X"b4388b19",
X"3370bf06",
X"71810652",
X"43557480",
X"2e80e838",
X"7b81bf06",
X"55748f24",
X"80dd389a",
X"19335574",
X"80d5389c",
X"19335574",
X"802e80cb",
X"38f31e70",
X"585e8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387c51",
X"ecf73f83",
X"e0800841",
X"83e08008",
X"8738901d",
X"08fea538",
X"80603475",
X"802e8838",
X"7d527f51",
X"83b13f60",
X"802e8638",
X"800b901e",
X"0c605660",
X"832e0981",
X"06883880",
X"0b901e0c",
X"85396081",
X"d238891f",
X"57901d08",
X"802e81a8",
X"38805675",
X"19703351",
X"5574a02e",
X"a0387485",
X"2e098106",
X"843881e5",
X"55747770",
X"81055934",
X"81167081",
X"ff065755",
X"877627d7",
X"38881933",
X"5574a02e",
X"a938ae77",
X"70810559",
X"34885675",
X"19703351",
X"5574a02e",
X"95387477",
X"70810559",
X"34811670",
X"81ff0657",
X"558a7627",
X"e2388b19",
X"337f8805",
X"349f1933",
X"9e1a3371",
X"982b7190",
X"2b079d1c",
X"3370882b",
X"72079c1e",
X"33710764",
X"0c52991d",
X"33981e33",
X"71882b07",
X"53515357",
X"5956747f",
X"84052397",
X"1933961a",
X"3371882b",
X"07565674",
X"7f860523",
X"8077347c",
X"51eafe3f",
X"83e08008",
X"5683e080",
X"08832e09",
X"81068838",
X"800b901e",
X"0c805696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"81b13f75",
X"83e0800c",
X"9e3d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"e0800c84",
X"3d0d04fc",
X"3d0d7655",
X"7483e680",
X"082eaf38",
X"80537451",
X"87cd3f83",
X"e0800881",
X"ff06ff14",
X"7081ff06",
X"7230709f",
X"2a515255",
X"53547280",
X"2e843871",
X"dd3873fe",
X"387483e6",
X"800c863d",
X"0d04ff3d",
X"0dff0b83",
X"e6800c84",
X"af3f8151",
X"87913f83",
X"e0800881",
X"ff065271",
X"ee3881d6",
X"3f7183e0",
X"800c833d",
X"0d04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"823f7280",
X"2ea03883",
X"e6941433",
X"75708105",
X"57348114",
X"7083ffff",
X"06ff1570",
X"83ffff06",
X"56525552",
X"dd39800b",
X"83e0800c",
X"863d0d04",
X"fc3d0d76",
X"787a1156",
X"53558053",
X"71742e93",
X"38721551",
X"703383e6",
X"94133481",
X"12811454",
X"52ea3980",
X"0b83e080",
X"0c863d0d",
X"04fd3d0d",
X"905483e6",
X"80085187",
X"803f83e0",
X"800881ff",
X"06ff1571",
X"30713070",
X"73079f2a",
X"729f2a06",
X"52555255",
X"5372db38",
X"853d0d04",
X"ff3d0d83",
X"e68c0810",
X"83e68408",
X"0780fce4",
X"0852710c",
X"833d0d04",
X"800b83e6",
X"8c0ce13f",
X"04810b83",
X"e68c0cd8",
X"3f04ed3f",
X"047183e6",
X"880c0480",
X"3d0d8051",
X"f43f810b",
X"83e68c0c",
X"810b83e6",
X"840cffb8",
X"3f823d0d",
X"04803d0d",
X"72307074",
X"07802583",
X"e6840c51",
X"ffa23f82",
X"3d0d04fe",
X"3d0d0293",
X"053380fc",
X"e8085473",
X"0c80fce4",
X"08527108",
X"70810651",
X"5170f738",
X"72087081",
X"ff0683e0",
X"800c5184",
X"3d0d0480",
X"3d0d81ff",
X"51cd3f83",
X"e0800881",
X"ff0683e0",
X"800c823d",
X"0d04ff3d",
X"0d74902b",
X"740780fc",
X"d8085271",
X"0c833d0d",
X"0404fb3d",
X"0d780284",
X"059f0533",
X"70982b55",
X"57557280",
X"259b3875",
X"80ff0656",
X"805280f7",
X"51e03f83",
X"e0800881",
X"ff065473",
X"812680ff",
X"388051fe",
X"e03fff9f",
X"3f8151fe",
X"d83fff97",
X"3f7551fe",
X"e63f7498",
X"2a51fedf",
X"3f74902a",
X"7081ff06",
X"5253fed3",
X"3f74882a",
X"7081ff06",
X"5253fec7",
X"3f7481ff",
X"0651febf",
X"3f815575",
X"80c02e09",
X"81068638",
X"8195558d",
X"397580c8",
X"2e098106",
X"84388187",
X"557451fe",
X"9e3f8a55",
X"fec53f83",
X"e0800881",
X"ff067098",
X"2b545472",
X"80258c38",
X"ff157081",
X"ff065653",
X"74e23873",
X"83e0800c",
X"873d0d04",
X"fa3d0dfd",
X"be3f8051",
X"fdd33f8a",
X"54fe903f",
X"ff147081",
X"ff065553",
X"73f33873",
X"74535580",
X"c051fea6",
X"3f83e080",
X"0881ff06",
X"5473812e",
X"09810682",
X"a13883aa",
X"5280c851",
X"fe8c3f83",
X"e0800881",
X"ff065372",
X"812e0981",
X"0681a938",
X"7454873d",
X"74115456",
X"fdc53f83",
X"e0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e538029a",
X"05335372",
X"812e0981",
X"0681db38",
X"029b0533",
X"5380ce90",
X"547281aa",
X"2e8e3881",
X"c93980e4",
X"51ff9fc0",
X"3fff1454",
X"73802e81",
X"b938820a",
X"5281e951",
X"fda43f83",
X"e0800881",
X"ff065372",
X"dd387252",
X"80fa51fd",
X"913f83e0",
X"800881ff",
X"06537281",
X"91387254",
X"731653fc",
X"d23f83e0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e8",
X"38873d33",
X"70862a70",
X"81065154",
X"548c5572",
X"80e43884",
X"5580df39",
X"745281e9",
X"51fccb3f",
X"83e08008",
X"81ff0653",
X"825581e9",
X"56817327",
X"86387355",
X"80c15680",
X"ce90548b",
X"3980e451",
X"ff9eb13f",
X"ff145473",
X"802ea938",
X"80527551",
X"fc983f83",
X"e0800881",
X"ff065372",
X"e0388480",
X"5280d051",
X"fc843f83",
X"e0800881",
X"ff065372",
X"802e8338",
X"80557483",
X"e6903480",
X"51fafe3f",
X"fbbd3f88",
X"3d0d04fb",
X"3d0d7754",
X"800b83e6",
X"90337083",
X"2a708106",
X"51555755",
X"72752e09",
X"81068538",
X"73892b54",
X"735280d1",
X"51fbbb3f",
X"83e08008",
X"81ff0653",
X"72bd3882",
X"b8c054fa",
X"fe3f83e0",
X"800881ff",
X"06537281",
X"ff2e0981",
X"068938ff",
X"145473e7",
X"389f3972",
X"81fe2e09",
X"81069638",
X"83ea9452",
X"83e69451",
X"fae83ffa",
X"ce3ffacb",
X"3f833981",
X"558051fa",
X"803ffabf",
X"3f7481ff",
X"0683e080",
X"0c873d0d",
X"04fb3d0d",
X"7783e694",
X"56548151",
X"f9e33f83",
X"e6903370",
X"832a7081",
X"06515456",
X"72853873",
X"892b5473",
X"5280d851",
X"fab43f83",
X"e0800881",
X"ff065372",
X"80e53881",
X"ff51f9cb",
X"3f81fe51",
X"f9c53f84",
X"80537470",
X"81055633",
X"51f9b83f",
X"ff137083",
X"ffff0651",
X"5372eb38",
X"7251f9a7",
X"3f7251f9",
X"a23ff9cb",
X"3f83e080",
X"089f0653",
X"a7885472",
X"852e8d38",
X"9a3980e4",
X"51ff9be8",
X"3fff1454",
X"f9ad3f83",
X"e0800881",
X"ff2e8438",
X"73e83880",
X"51f8da3f",
X"f9993f80",
X"0b83e080",
X"0c873d0d",
X"0483e08c",
X"080283e0",
X"8c0cfd3d",
X"0d805383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"05085183",
X"d43f83e0",
X"80087083",
X"e0800c54",
X"853d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cfd3d0d",
X"815383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"085183a1",
X"3f83e080",
X"087083e0",
X"800c5485",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"f93d0d80",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"88050880",
X"25b93883",
X"e08c0888",
X"05083083",
X"e08c0888",
X"050c800b",
X"83e08c08",
X"f4050c83",
X"e08c08fc",
X"05088a38",
X"810b83e0",
X"8c08f405",
X"0c83e08c",
X"08f40508",
X"83e08c08",
X"fc050c83",
X"e08c088c",
X"05088025",
X"b93883e0",
X"8c088c05",
X"083083e0",
X"8c088c05",
X"0c800b83",
X"e08c08f0",
X"050c83e0",
X"8c08fc05",
X"088a3881",
X"0b83e08c",
X"08f0050c",
X"83e08c08",
X"f0050883",
X"e08c08fc",
X"050c8053",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"81df3f83",
X"e0800870",
X"83e08c08",
X"f8050c54",
X"83e08c08",
X"fc050880",
X"2e903883",
X"e08c08f8",
X"05083083",
X"e08c08f8",
X"050c83e0",
X"8c08f805",
X"087083e0",
X"800c5489",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"fb3d0d80",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"88050880",
X"25993883",
X"e08c0888",
X"05083083",
X"e08c0888",
X"050c810b",
X"83e08c08",
X"fc050c83",
X"e08c088c",
X"05088025",
X"903883e0",
X"8c088c05",
X"083083e0",
X"8c088c05",
X"0c815383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"050851bd",
X"3f83e080",
X"087083e0",
X"8c08f805",
X"0c5483e0",
X"8c08fc05",
X"08802e90",
X"3883e08c",
X"08f80508",
X"3083e08c",
X"08f8050c",
X"83e08c08",
X"f8050870",
X"83e0800c",
X"54873d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cfd3d",
X"0d810b83",
X"e08c08fc",
X"050c800b",
X"83e08c08",
X"f8050c83",
X"e08c088c",
X"050883e0",
X"8c088805",
X"0827b938",
X"83e08c08",
X"fc050880",
X"2eae3880",
X"0b83e08c",
X"088c0508",
X"24a23883",
X"e08c088c",
X"05081083",
X"e08c088c",
X"050c83e0",
X"8c08fc05",
X"081083e0",
X"8c08fc05",
X"0cffb839",
X"83e08c08",
X"fc050880",
X"2e80e138",
X"83e08c08",
X"8c050883",
X"e08c0888",
X"050826ad",
X"3883e08c",
X"08880508",
X"83e08c08",
X"8c050831",
X"83e08c08",
X"88050c83",
X"e08c08f8",
X"050883e0",
X"8c08fc05",
X"080783e0",
X"8c08f805",
X"0c83e08c",
X"08fc0508",
X"812a83e0",
X"8c08fc05",
X"0c83e08c",
X"088c0508",
X"812a83e0",
X"8c088c05",
X"0cff9539",
X"83e08c08",
X"90050880",
X"2e933883",
X"e08c0888",
X"05087083",
X"e08c08f4",
X"050c5191",
X"3983e08c",
X"08f80508",
X"7083e08c",
X"08f4050c",
X"5183e08c",
X"08f40508",
X"83e0800c",
X"853d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cff3d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"8106ff11",
X"70097083",
X"e08c088c",
X"05080683",
X"e08c08fc",
X"05081183",
X"e08c08fc",
X"050c83e0",
X"8c088805",
X"08812a83",
X"e08c0888",
X"050c83e0",
X"8c088c05",
X"081083e0",
X"8c088c05",
X"0c515151",
X"5183e08c",
X"08880508",
X"802e8438",
X"ffab3983",
X"e08c08fc",
X"05087083",
X"e0800c51",
X"833d0d83",
X"e08c0c04",
X"fc3d0d76",
X"70797b55",
X"5555558f",
X"72278c38",
X"72750783",
X"06517080",
X"2ea938ff",
X"125271ff",
X"2e983872",
X"70810554",
X"33747081",
X"055634ff",
X"125271ff",
X"2e098106",
X"ea387483",
X"e0800c86",
X"3d0d0474",
X"51727084",
X"05540871",
X"70840553",
X"0c727084",
X"05540871",
X"70840553",
X"0c727084",
X"05540871",
X"70840553",
X"0c727084",
X"05540871",
X"70840553",
X"0cf01252",
X"718f26c9",
X"38837227",
X"95387270",
X"84055408",
X"71708405",
X"530cfc12",
X"52718326",
X"ed387054",
X"ff813900",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"000009a5",
X"000009e6",
X"00000a08",
X"00000a26",
X"00000a26",
X"00000a26",
X"00000a26",
X"00000a95",
X"00000ac5",
X"70704740",
X"9c704268",
X"9c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"43617274",
X"72696467",
X"6520386b",
X"2073696d",
X"706c6500",
X"45786974",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"25732025",
X"73000000",
X"2e2e0000",
X"2f000000",
X"41545200",
X"58464400",
X"58455800",
X"524f4d00",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"6e616d65",
X"20000000",
X"25303278",
X"00000000",
X"00000000",
X"00000000",
X"00003cb8",
X"00003cbc",
X"00003cc4",
X"00003cd0",
X"00003cdc",
X"00003ce8",
X"00003cf4",
X"00003cf8",
X"0001d20f",
X"0001d400",
X"0001d401",
X"0001d409",
X"0001d010",
X"0001d301",
X"0001d300",
X"0001d20a",
X"0001d01b",
X"0001d016",
X"0001d019",
X"0001d018",
X"0001d017",
X"0001d01a",
X"0001d403",
X"0001d402",
X"0001d40e",
X"0004007c",
X"00040078",
X"00040074",
X"00040068",
X"00040060",
X"0004005c",
X"00040058",
X"00040054",
X"00040050",
X"0004004c",
X"00040048",
X"00040044",
X"00040040",
X"00040034",
X"00040030",
X"0004002c",
X"00040028",
X"00040024",
X"00040020",
X"0004001c",
X"00040018",
X"00040014",
X"00040010",
X"0004000c",
X"00040008",
X"00040004",
X"00040000",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
