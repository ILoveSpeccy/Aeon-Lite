library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

entity chram is
   Port (
      CLK         : in  std_logic;
      CHRAM_A     : in  std_logic_vector(9 downto 0);
      CHRAM_WR    : in  std_logic;
      CHRAM_DI    : in  std_logic_vector(8 downto 0);
      CHRAM_DO    : out std_logic_vector(8 downto 0);
      CHRAM_VA    : in  std_logic_vector(9 downto 0);
      CHRAM_VD    : out std_logic_vector(8 downto 0)
   );
end chram;

architecture rtl of chram is

   subtype word_t is std_logic_vector(8 downto 0);
   type memory_t is array(0 to 1023) of word_t;
   shared variable ram : memory_t := (
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "001000011", "001010000", "000101111", "001001101", "000101101", "000111000", "000110000", "000100000", 
      "000100000", "001110110", "000101110", "000100000", "000110010", "000101110", "000110010", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "011101111", "011100110", "011110000", "000100000", "000100000", "011101110", "011101001", "011101001", 
      "011110001", "011100110", "000100000", "000100000", "011101101", "011100111", "011110101", "000100000", 
      "000100000", "001000010", "001001001", "001001111", "001010011", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "001010110", "001100101", "001110010", "000101110", "000100000", "000110001", "000101110", "000110010", 
      "000100000", "000101000", "001100011", "000101001", "000100000", "001001001", "001001001", "001001001", 
      "000100000", "000110001", "000111001", "000111000", "000111000", "000100000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "001000001", "000111110", "001000100", "001001001", "001010010", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "001000001", "000111010", "000100000", "001000010", "001001001", "001001110", "001000001", "001001100", 
      "001000101", "001001110", "001000100", "000100000", "001000011", "001001111", "001001101", "000100000", 
      "000111010", "000100000", "001000011", "001001000", "001000001", "001010011", "001000101", "001010010", 
      "000100000", "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", "000111010", 
      "000100000", "001001010", "001000001", "001001101", "001010000", "001000101", "001010010", "000100000", 
      "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", "000111010", "000100000", 
      "001001011", "001001100", "001000001", "001000100", "000110001", "000100000", "000100000", "000100000", 
      "000100000", "001000011", "001001111", "001001101", "000000000", "000000000", "000000000", "000000000", 
      "001000001", "000111010", "000100000", "001001101", "001000001", "001000110", "001001001", "001000001", 
      "000100000", "000100000", "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", 
      "000111010", "000100000", "001010000", "001000001", "001000011", "001001101", "001000001", "001001110", 
      "000100000", "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", "000111010", 
      "000100000", "001010000", "001001111", "001010000", "001001011", "001001111", "001010010", "001001110", 
      "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", "000111010", "000100000", 
      "001010011", "001001111", "001001011", "001001111", "000100000", "000100000", "000100000", "000100000", 
      "000100000", "001000011", "001001111", "001001101", "000000000", "000000000", "000000000", "000000000", 
      "001000001", "000111010", "000100000", "001010011", "001010100", "001000001", "001001100", "001001011", 
      "001000101", "001010010", "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", 
      "000111010", "000100000", "001011000", "001011001", "001011010", "001001111", "001001110", "000100000", 
      "000100000", "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", "000111010", 
      "000100000", "001011010", "001010111", "000100000", "000100000", "000100000", "000100000", "000100000", 
      "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", "000111010", "000100000", 
      "001000110", "001000001", "001001001", "001010010", "000100000", "000100000", "000100000", "000100000", 
      "000100000", "001000011", "001001111", "001001101", "000000000", "000000000", "000000000", "000000000", 
      "001000001", "000111010", "000100000", "001000010", "001001111", "001001101", "001000010", "001000101", 
      "001010010", "000100000", "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", 
      "000111010", "000100000", "001000011", "001001111", "001001100", "001001111", "001010010", "001000010", 
      "001000001", "001001100", "000100000", "001000011", "001001111", "001001101", "000100000", "000111010", 
      "000100000", "001000110", "001001001", "001010110", "001010100", "001000101", "001000101", "001001110", 
      "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", "000111010", "000100000", 
      "001010011", "001000001", "001001101", "001001111", "001010110", "001000001", "001010010", "000100000", 
      "000100000", "001000011", "001001111", "001001101", "000000000", "000000000", "000000000", "000000000", 
      "001000001", "000111010", "000100000", "001011000", "001000001", "001010010", "001010100", "000100000", 
      "000100000", "000100000", "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", 
      "000111010", "000100000", "001000001", "001001110", "001010100", "001001111", "001001110", "000100000", 
      "000100000", "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", "000111010", 
      "000100000", "001010010", "001000001", "001001100", "001001100", "001011001", "000100000", "000100000", 
      "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", "000111010", "000100000", 
      "001010100", "001000101", "001010100", "001010010", "001001001", "001010011", "000100000", "000100000", 
      "000100000", "001000011", "001001111", "001001101", "000000000", "000000000", "000000000", "000000000", 
      "001000001", "000111010", "000100000", "001000010", "001000001", "001010010", "001010011", "000100000", 
      "000100000", "000100000", "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", 
      "000111010", "000100000", "001000011", "001001001", "001010010", "001000011", "001010101", "001010011", 
      "000100000", "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", "000111010", 
      "000100000", "001000011", "001001001", "001010010", "001000011", "001010101", "001010011", "000100000", 
      "000100000", "000100000", "001000100", "001000001", "001010100", "000100000", "000111010", "000100000", 
      "001000011", "001001001", "001010010", "001000011", "001010101", "001010011", "000100000", "000100000", 
      "000100000", "001010000", "001000011", "000110001", "000000000", "000000000", "000000000", "000000000", 
      "001000001", "000111010", "000100000", "001000011", "001001001", "001010010", "001000011", "001010101", 
      "001010011", "000110000", "000100000", "000100000", "001010010", "001000101", "001011010", "000100000", 
      "000111010", "000100000", "001000011", "001001001", "001010010", "001000011", "001010101", "001010011", 
      "000110001", "000100000", "000100000", "001010010", "001000101", "001011010", "000100000", "000111010", 
      "000100000", "001000011", "001001001", "001010010", "001000011", "001010101", "001010011", "000110100", 
      "000100000", "000100000", "001010010", "001000101", "001011010", "000100000", "000111010", "000100000", 
      "001000011", "001001001", "001010010", "001000011", "001010101", "001010011", "000110101", "000100000", 
      "000100000", "001010010", "001000101", "001011010", "000000000", "000000000", "000000000", "000000000", 
      "001000001", "000111010", "000100000", "001000011", "001001001", "001010010", "001000011", "001010101", 
      "001010011", "000111001", "000100000", "000100000", "001010010", "001000101", "001011010", "000100000", 
      "000111010", "000100000", "001010000", "001000001", "001000111", "001000001", "001001110", "001001001", 
      "001001110", "001001001", "000100000", "001000011", "001001111", "001001101", "000100000", "000111010", 
      "000100000", "001010011", "001010000", "001001111", "001010010", "001010100", "000100000", "000100000", 
      "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", "000111010", "000100000", 
      "001000111", "001000001", "001001100", "001000001", "001011000", "001001001", "001000001", "001001110", 
      "000100000", "001000011", "001001111", "001001101", "000000000", "000000000", "000000000", "000000000", 
      "001000001", "000111010", "000100000", "001010011", "001001111", "001001111", "000100000", "000100000", 
      "000100000", "000100000", "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", 
      "000111010", "000100000", "001001110", "001001001", "001001110", "001001010", "001000001", "000100000", 
      "000100000", "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", "000111010", 
      "000100000", "001001011", "000110010", "000100000", "000100000", "000100000", "000100000", "000100000", 
      "000100000", "000100000", "001000011", "001001111", "001001101", "000100000", "000111010", "000100000", 
      "001010100", "001010010", "001000101", "001000001", "001010011", "000100000", "000100000", "000100000", 
      "000100000", "001000011", "001001111", "001001101", "000000000", "000000000", "000000000", "000000000", 
      "001000001", "000111110", "100000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", 
      "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000" );

begin

   process(CLK)
   begin
      if rising_edge(CLK) then 
         if CHRAM_WR = '1' then
            ram(to_integer(unsigned(CHRAM_A))) := CHRAM_DI;
         else
            CHRAM_DO <= ram(to_integer(unsigned(CHRAM_A)));
         end if;
      end if;
   end process;   
   
   process(CLK)
   begin
      if rising_edge(CLK) then 
         CHRAM_VD <= ram(to_integer(unsigned(CHRAM_VA)));
      end if;
   end process;
 
end rtl;
