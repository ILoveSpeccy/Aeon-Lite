---------------------------------------------------------------------------
-- (c) 2013 mark watson
-- I am happy for anyone to use this for non-commercial use.
-- If my vhdl files are used commercially or otherwise sold,
-- please contact me for explicit permission at scrameta (gmail).
-- This applies for source and binary form and derived works.
---------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use IEEE.STD_LOGIC_MISC.all;

ENTITY pokey_mixer IS
PORT 
( 
	CLK : IN STD_LOGIC;
	
	CHANNEL_ENABLE : IN STD_LOGIC_VECTOR(3 downto 0);
		
	CHANNEL_0 : IN STD_LOGIC_VECTOR(3 downto 0);
	CHANNEL_1 : IN STD_LOGIC_VECTOR(3 downto 0);
	CHANNEL_2 : IN STD_LOGIC_VECTOR(3 downto 0);
	CHANNEL_3 : IN STD_LOGIC_VECTOR(3 downto 0);
	
	GTIA_SOUND : IN STD_LOGIC;

	COVOX_CHANNEL_0 : IN STD_LOGIC_VECTOR(7 downto 0);
	COVOX_CHANNEL_1 : IN STD_LOGIC_VECTOR(7 downto 0);
	
	VOLUME_OUT : OUT STD_LOGIC_vector(15 downto 0)
);
END pokey_mixer;

ARCHITECTURE vhdl OF pokey_mixer IS
	signal volume_next : std_logic_vector(15 downto 0);
	signal volume_reg : std_logic_vector(15 downto 0);
	
	signal volume_sum : std_logic_vector(9 downto 0);
	
	signal channel_0_en : std_logic_vector(3 downto 0);
	signal channel_1_en : std_logic_vector(3 downto 0);
	signal channel_2_en : std_logic_vector(3 downto 0);
	signal channel_3_en : std_logic_vector(3 downto 0);
BEGIN
	-- register
	process(clk)
	begin
		if (clk'event and clk='1') then
			volume_reg <= volume_next;
		end if;
	end process;
	
	-- next state
	process(channel_enable,channel_0,channel_1,channel_2,channel_3)
	begin
		channel_0_en <= channel_0;
		channel_1_en <= channel_1;
		channel_2_en <= channel_2;
		channel_3_en <= channel_3;
	
--		if (channel_enable(3)='0') then
--			channel_0_en <= X"0";
--		end if;
--		
--		if (channel_enable(2)='0') then
--			channel_1_en <= X"0";
--		end if;
--
--		if (channel_enable(1)='0') then
--			channel_2_en <= X"0";
--		end if;
--		
--		if (channel_enable(0)='0') then
--			channel_3_en <= X"0";
--		end if;
	end process;
	
	process (channel_0_en,channel_1_en,channel_2_en,channel_3_en,covox_CHANNEL_0,covox_channel_1,gtia_sound)
		variable channel0_en_long : unsigned(10 downto 0);
		variable channel1_en_long : unsigned(10 downto 0);
		variable channel2_en_long : unsigned(10 downto 0);
		variable channel3_en_long : unsigned(10 downto 0);
		variable gtia_sound_long : unsigned(10 downto 0);
		variable covox_0_long : unsigned(10 downto 0);
		variable covox_1_long : unsigned(10 downto 0);
		
		variable volume_int_sum : unsigned(10 downto 0);
	begin
		channel0_en_long := (others=>'0');
		channel1_en_long := (others=>'0');
		channel2_en_long := (others=>'0');
		channel3_en_long := (others=>'0');
		gtia_sound_long := (others=>'0');
		covox_0_long := (others=>'0');
		covox_1_long := (others=>'0');

		channel0_en_long(7 downto 4) := unsigned(channel_0_en);
		channel1_en_long(7 downto 4) := unsigned(channel_1_en);
		channel2_en_long(7 downto 4) := unsigned(channel_2_en);
		channel3_en_long(7 downto 4) := unsigned(channel_3_en);
		gtia_sound_long(7 downto 4) := gtia_sound&gtia_sound&gtia_sound&gtia_sound;
		covox_0_long(7 downto 0) := unsigned(covox_channel_0);
		covox_1_long(7 downto 0) := unsigned(covox_channel_1);

		volume_int_sum := ((channel0_en_long + channel1_en_long) + (channel2_en_long + channel3_en_long)) + (gtia_sound_long + (covox_0_long + covox_1_long));

		volume_sum(8 downto 0) <= std_logic_vector(volume_int_sum(8 downto 0));
		volume_sum(9) <= volume_int_sum(10) or volume_int_sum(9);
	end process;
	
 	process (volume_sum, volume_next)
	begin
		case volume_sum(9 downto 0) is 
			when "0000000000" =>
				volume_next <= X"0000";
			when "0000000001" =>
				volume_next <= X"00cc";
			when "0000000010" =>
				volume_next <= X"0198";
			when "0000000011" =>
				volume_next <= X"0264";
			when "0000000100" =>
				volume_next <= X"032f";
			when "0000000101" =>
				volume_next <= X"03fa";
			when "0000000110" =>
				volume_next <= X"04c4";
			when "0000000111" =>
				volume_next <= X"058e";
			when "0000001000" =>
				volume_next <= X"0657";
			when "0000001001" =>
				volume_next <= X"0720";
			when "0000001010" =>
				volume_next <= X"07e8";
			when "0000001011" =>
				volume_next <= X"08b0";
			when "0000001100" =>
				volume_next <= X"0977";
			when "0000001101" =>
				volume_next <= X"0a3e";
			when "0000001110" =>
				volume_next <= X"0b05";
			when "0000001111" =>
				volume_next <= X"0bcb";
			when "0000010000" =>
				volume_next <= X"0c91";
			when "0000010001" =>
				volume_next <= X"0d56";
			when "0000010010" =>
				volume_next <= X"0e1a";
			when "0000010011" =>
				volume_next <= X"0edf";
			when "0000010100" =>
				volume_next <= X"0fa2";
			when "0000010101" =>
				volume_next <= X"1066";
			when "0000010110" =>
				volume_next <= X"1128";
			when "0000010111" =>
				volume_next <= X"11eb";
			when "0000011000" =>
				volume_next <= X"12ad";
			when "0000011001" =>
				volume_next <= X"136e";
			when "0000011010" =>
				volume_next <= X"142f";
			when "0000011011" =>
				volume_next <= X"14f0";
			when "0000011100" =>
				volume_next <= X"15b0";
			when "0000011101" =>
				volume_next <= X"1670";
			when "0000011110" =>
				volume_next <= X"172f";
			when "0000011111" =>
				volume_next <= X"17ee";
			when "0000100000" =>
				volume_next <= X"18ac";
			when "0000100001" =>
				volume_next <= X"196a";
			when "0000100010" =>
				volume_next <= X"1a27";
			when "0000100011" =>
				volume_next <= X"1ae4";
			when "0000100100" =>
				volume_next <= X"1ba1";
			when "0000100101" =>
				volume_next <= X"1c5d";
			when "0000100110" =>
				volume_next <= X"1d18";
			when "0000100111" =>
				volume_next <= X"1dd3";
			when "0000101000" =>
				volume_next <= X"1e8e";
			when "0000101001" =>
				volume_next <= X"1f48";
			when "0000101010" =>
				volume_next <= X"2002";
			when "0000101011" =>
				volume_next <= X"20bc";
			when "0000101100" =>
				volume_next <= X"2174";
			when "0000101101" =>
				volume_next <= X"222d";
			when "0000101110" =>
				volume_next <= X"22e5";
			when "0000101111" =>
				volume_next <= X"239d";
			when "0000110000" =>
				volume_next <= X"2454";
			when "0000110001" =>
				volume_next <= X"250a";
			when "0000110010" =>
				volume_next <= X"25c1";
			when "0000110011" =>
				volume_next <= X"2677";
			when "0000110100" =>
				volume_next <= X"272c";
			when "0000110101" =>
				volume_next <= X"27e1";
			when "0000110110" =>
				volume_next <= X"2895";
			when "0000110111" =>
				volume_next <= X"2949";
			when "0000111000" =>
				volume_next <= X"29fd";
			when "0000111001" =>
				volume_next <= X"2ab0";
			when "0000111010" =>
				volume_next <= X"2b63";
			when "0000111011" =>
				volume_next <= X"2c15";
			when "0000111100" =>
				volume_next <= X"2cc7";
			when "0000111101" =>
				volume_next <= X"2d79";
			when "0000111110" =>
				volume_next <= X"2e2a";
			when "0000111111" =>
				volume_next <= X"2eda";
			when "0001000000" =>
				volume_next <= X"2f8b";
			when "0001000001" =>
				volume_next <= X"303a";
			when "0001000010" =>
				volume_next <= X"30ea";
			when "0001000011" =>
				volume_next <= X"3198";
			when "0001000100" =>
				volume_next <= X"3247";
			when "0001000101" =>
				volume_next <= X"32f5";
			when "0001000110" =>
				volume_next <= X"33a2";
			when "0001000111" =>
				volume_next <= X"3450";
			when "0001001000" =>
				volume_next <= X"34fc";
			when "0001001001" =>
				volume_next <= X"35a9";
			when "0001001010" =>
				volume_next <= X"3654";
			when "0001001011" =>
				volume_next <= X"3700";
			when "0001001100" =>
				volume_next <= X"37ab";
			when "0001001101" =>
				volume_next <= X"3856";
			when "0001001110" =>
				volume_next <= X"3900";
			when "0001001111" =>
				volume_next <= X"39a9";
			when "0001010000" =>
				volume_next <= X"3a53";
			when "0001010001" =>
				volume_next <= X"3afc";
			when "0001010010" =>
				volume_next <= X"3ba4";
			when "0001010011" =>
				volume_next <= X"3c4c";
			when "0001010100" =>
				volume_next <= X"3cf4";
			when "0001010101" =>
				volume_next <= X"3d9b";
			when "0001010110" =>
				volume_next <= X"3e42";
			when "0001010111" =>
				volume_next <= X"3ee8";
			when "0001011000" =>
				volume_next <= X"3f8e";
			when "0001011001" =>
				volume_next <= X"4034";
			when "0001011010" =>
				volume_next <= X"40d9";
			when "0001011011" =>
				volume_next <= X"417d";
			when "0001011100" =>
				volume_next <= X"4222";
			when "0001011101" =>
				volume_next <= X"42c5";
			when "0001011110" =>
				volume_next <= X"4369";
			when "0001011111" =>
				volume_next <= X"440c";
			when "0001100000" =>
				volume_next <= X"44af";
			when "0001100001" =>
				volume_next <= X"4551";
			when "0001100010" =>
				volume_next <= X"45f3";
			when "0001100011" =>
				volume_next <= X"4694";
			when "0001100100" =>
				volume_next <= X"4735";
			when "0001100101" =>
				volume_next <= X"47d5";
			when "0001100110" =>
				volume_next <= X"4876";
			when "0001100111" =>
				volume_next <= X"4915";
			when "0001101000" =>
				volume_next <= X"49b5";
			when "0001101001" =>
				volume_next <= X"4a53";
			when "0001101010" =>
				volume_next <= X"4af2";
			when "0001101011" =>
				volume_next <= X"4b90";
			when "0001101100" =>
				volume_next <= X"4c2e";
			when "0001101101" =>
				volume_next <= X"4ccb";
			when "0001101110" =>
				volume_next <= X"4d68";
			when "0001101111" =>
				volume_next <= X"4e04";
			when "0001110000" =>
				volume_next <= X"4ea0";
			when "0001110001" =>
				volume_next <= X"4f3c";
			when "0001110010" =>
				volume_next <= X"4fd7";
			when "0001110011" =>
				volume_next <= X"5072";
			when "0001110100" =>
				volume_next <= X"510d";
			when "0001110101" =>
				volume_next <= X"51a7";
			when "0001110110" =>
				volume_next <= X"5240";
			when "0001110111" =>
				volume_next <= X"52da";
			when "0001111000" =>
				volume_next <= X"5372";
			when "0001111001" =>
				volume_next <= X"540b";
			when "0001111010" =>
				volume_next <= X"54a3";
			when "0001111011" =>
				volume_next <= X"553a";
			when "0001111100" =>
				volume_next <= X"55d2";
			when "0001111101" =>
				volume_next <= X"5669";
			when "0001111110" =>
				volume_next <= X"56ff";
			when "0001111111" =>
				volume_next <= X"5795";
			when "0010000000" =>
				volume_next <= X"582b";
			when "0010000001" =>
				volume_next <= X"58c0";
			when "0010000010" =>
				volume_next <= X"5955";
			when "0010000011" =>
				volume_next <= X"59e9";
			when "0010000100" =>
				volume_next <= X"5a7d";
			when "0010000101" =>
				volume_next <= X"5b11";
			when "0010000110" =>
				volume_next <= X"5ba4";
			when "0010000111" =>
				volume_next <= X"5c37";
			when "0010001000" =>
				volume_next <= X"5cca";
			when "0010001001" =>
				volume_next <= X"5d5c";
			when "0010001010" =>
				volume_next <= X"5dee";
			when "0010001011" =>
				volume_next <= X"5e7f";
			when "0010001100" =>
				volume_next <= X"5f10";
			when "0010001101" =>
				volume_next <= X"5fa0";
			when "0010001110" =>
				volume_next <= X"6031";
			when "0010001111" =>
				volume_next <= X"60c0";
			when "0010010000" =>
				volume_next <= X"6150";
			when "0010010001" =>
				volume_next <= X"61df";
			when "0010010010" =>
				volume_next <= X"626d";
			when "0010010011" =>
				volume_next <= X"62fc";
			when "0010010100" =>
				volume_next <= X"638a";
			when "0010010101" =>
				volume_next <= X"6417";
			when "0010010110" =>
				volume_next <= X"64a4";
			when "0010010111" =>
				volume_next <= X"6531";
			when "0010011000" =>
				volume_next <= X"65bd";
			when "0010011001" =>
				volume_next <= X"6649";
			when "0010011010" =>
				volume_next <= X"66d5";
			when "0010011011" =>
				volume_next <= X"6760";
			when "0010011100" =>
				volume_next <= X"67eb";
			when "0010011101" =>
				volume_next <= X"6875";
			when "0010011110" =>
				volume_next <= X"68ff";
			when "0010011111" =>
				volume_next <= X"6989";
			when "0010100000" =>
				volume_next <= X"6a12";
			when "0010100001" =>
				volume_next <= X"6a9b";
			when "0010100010" =>
				volume_next <= X"6b23";
			when "0010100011" =>
				volume_next <= X"6bac";
			when "0010100100" =>
				volume_next <= X"6c33";
			when "0010100101" =>
				volume_next <= X"6cbb";
			when "0010100110" =>
				volume_next <= X"6d42";
			when "0010100111" =>
				volume_next <= X"6dc9";
			when "0010101000" =>
				volume_next <= X"6e4f";
			when "0010101001" =>
				volume_next <= X"6ed5";
			when "0010101010" =>
				volume_next <= X"6f5a";
			when "0010101011" =>
				volume_next <= X"6fdf";
			when "0010101100" =>
				volume_next <= X"7064";
			when "0010101101" =>
				volume_next <= X"70e9";
			when "0010101110" =>
				volume_next <= X"716d";
			when "0010101111" =>
				volume_next <= X"71f0";
			when "0010110000" =>
				volume_next <= X"7274";
			when "0010110001" =>
				volume_next <= X"72f7";
			when "0010110010" =>
				volume_next <= X"7379";
			when "0010110011" =>
				volume_next <= X"73fc";
			when "0010110100" =>
				volume_next <= X"747d";
			when "0010110101" =>
				volume_next <= X"74ff";
			when "0010110110" =>
				volume_next <= X"7580";
			when "0010110111" =>
				volume_next <= X"7601";
			when "0010111000" =>
				volume_next <= X"7681";
			when "0010111001" =>
				volume_next <= X"7701";
			when "0010111010" =>
				volume_next <= X"7781";
			when "0010111011" =>
				volume_next <= X"7800";
			when "0010111100" =>
				volume_next <= X"787f";
			when "0010111101" =>
				volume_next <= X"78fe";
			when "0010111110" =>
				volume_next <= X"797c";
			when "0010111111" =>
				volume_next <= X"79fa";
			when "0011000000" =>
				volume_next <= X"7a77";
			when "0011000001" =>
				volume_next <= X"7af5";
			when "0011000010" =>
				volume_next <= X"7b71";
			when "0011000011" =>
				volume_next <= X"7bee";
			when "0011000100" =>
				volume_next <= X"7c6a";
			when "0011000101" =>
				volume_next <= X"7ce6";
			when "0011000110" =>
				volume_next <= X"7d61";
			when "0011000111" =>
				volume_next <= X"7ddc";
			when "0011001000" =>
				volume_next <= X"7e57";
			when "0011001001" =>
				volume_next <= X"7ed1";
			when "0011001010" =>
				volume_next <= X"7f4b";
			when "0011001011" =>
				volume_next <= X"7fc5";
			when "0011001100" =>
				volume_next <= X"803e";
			when "0011001101" =>
				volume_next <= X"80b7";
			when "0011001110" =>
				volume_next <= X"812f";
			when "0011001111" =>
				volume_next <= X"81a7";
			when "0011010000" =>
				volume_next <= X"821f";
			when "0011010001" =>
				volume_next <= X"8297";
			when "0011010010" =>
				volume_next <= X"830e";
			when "0011010011" =>
				volume_next <= X"8385";
			when "0011010100" =>
				volume_next <= X"83fb";
			when "0011010101" =>
				volume_next <= X"8471";
			when "0011010110" =>
				volume_next <= X"84e7";
			when "0011010111" =>
				volume_next <= X"855d";
			when "0011011000" =>
				volume_next <= X"85d2";
			when "0011011001" =>
				volume_next <= X"8646";
			when "0011011010" =>
				volume_next <= X"86bb";
			when "0011011011" =>
				volume_next <= X"872f";
			when "0011011100" =>
				volume_next <= X"87a2";
			when "0011011101" =>
				volume_next <= X"8816";
			when "0011011110" =>
				volume_next <= X"8889";
			when "0011011111" =>
				volume_next <= X"88fc";
			when "0011100000" =>
				volume_next <= X"896e";
			when "0011100001" =>
				volume_next <= X"89e0";
			when "0011100010" =>
				volume_next <= X"8a51";
			when "0011100011" =>
				volume_next <= X"8ac3";
			when "0011100100" =>
				volume_next <= X"8b34";
			when "0011100101" =>
				volume_next <= X"8ba4";
			when "0011100110" =>
				volume_next <= X"8c15";
			when "0011100111" =>
				volume_next <= X"8c85";
			when "0011101000" =>
				volume_next <= X"8cf4";
			when "0011101001" =>
				volume_next <= X"8d64";
			when "0011101010" =>
				volume_next <= X"8dd3";
			when "0011101011" =>
				volume_next <= X"8e41";
			when "0011101100" =>
				volume_next <= X"8eaf";
			when "0011101101" =>
				volume_next <= X"8f1d";
			when "0011101110" =>
				volume_next <= X"8f8b";
			when "0011101111" =>
				volume_next <= X"8ff8";
			when "0011110000" =>
				volume_next <= X"9065";
			when "0011110001" =>
				volume_next <= X"90d2";
			when "0011110010" =>
				volume_next <= X"913e";
			when "0011110011" =>
				volume_next <= X"91aa";
			when "0011110100" =>
				volume_next <= X"9216";
			when "0011110101" =>
				volume_next <= X"9281";
			when "0011110110" =>
				volume_next <= X"92ec";
			when "0011110111" =>
				volume_next <= X"9357";
			when "0011111000" =>
				volume_next <= X"93c1";
			when "0011111001" =>
				volume_next <= X"942b";
			when "0011111010" =>
				volume_next <= X"9495";
			when "0011111011" =>
				volume_next <= X"94fe";
			when "0011111100" =>
				volume_next <= X"9567";
			when "0011111101" =>
				volume_next <= X"95d0";
			when "0011111110" =>
				volume_next <= X"9638";
			when "0011111111" =>
				volume_next <= X"96a0";
			when "0100000000" =>
				volume_next <= X"9708";
			when "0100000001" =>
				volume_next <= X"9770";
			when "0100000010" =>
				volume_next <= X"97d7";
			when "0100000011" =>
				volume_next <= X"983d";
			when "0100000100" =>
				volume_next <= X"98a4";
			when "0100000101" =>
				volume_next <= X"990a";
			when "0100000110" =>
				volume_next <= X"9970";
			when "0100000111" =>
				volume_next <= X"99d5";
			when "0100001000" =>
				volume_next <= X"9a3b";
			when "0100001001" =>
				volume_next <= X"9a9f";
			when "0100001010" =>
				volume_next <= X"9b04";
			when "0100001011" =>
				volume_next <= X"9b68";
			when "0100001100" =>
				volume_next <= X"9bcc";
			when "0100001101" =>
				volume_next <= X"9c30";
			when "0100001110" =>
				volume_next <= X"9c93";
			when "0100001111" =>
				volume_next <= X"9cf6";
			when "0100010000" =>
				volume_next <= X"9d59";
			when "0100010001" =>
				volume_next <= X"9dbb";
			when "0100010010" =>
				volume_next <= X"9e1d";
			when "0100010011" =>
				volume_next <= X"9e7f";
			when "0100010100" =>
				volume_next <= X"9ee0";
			when "0100010101" =>
				volume_next <= X"9f41";
			when "0100010110" =>
				volume_next <= X"9fa2";
			when "0100010111" =>
				volume_next <= X"a003";
			when "0100011000" =>
				volume_next <= X"a063";
			when "0100011001" =>
				volume_next <= X"a0c3";
			when "0100011010" =>
				volume_next <= X"a122";
			when "0100011011" =>
				volume_next <= X"a182";
			when "0100011100" =>
				volume_next <= X"a1e1";
			when "0100011101" =>
				volume_next <= X"a23f";
			when "0100011110" =>
				volume_next <= X"a29e";
			when "0100011111" =>
				volume_next <= X"a2fc";
			when "0100100000" =>
				volume_next <= X"a359";
			when "0100100001" =>
				volume_next <= X"a3b7";
			when "0100100010" =>
				volume_next <= X"a414";
			when "0100100011" =>
				volume_next <= X"a471";
			when "0100100100" =>
				volume_next <= X"a4cd";
			when "0100100101" =>
				volume_next <= X"a52a";
			when "0100100110" =>
				volume_next <= X"a586";
			when "0100100111" =>
				volume_next <= X"a5e1";
			when "0100101000" =>
				volume_next <= X"a63c";
			when "0100101001" =>
				volume_next <= X"a698";
			when "0100101010" =>
				volume_next <= X"a6f2";
			when "0100101011" =>
				volume_next <= X"a74d";
			when "0100101100" =>
				volume_next <= X"a7a7";
			when "0100101101" =>
				volume_next <= X"a801";
			when "0100101110" =>
				volume_next <= X"a85a";
			when "0100101111" =>
				volume_next <= X"a8b4";
			when "0100110000" =>
				volume_next <= X"a90c";
			when "0100110001" =>
				volume_next <= X"a965";
			when "0100110010" =>
				volume_next <= X"a9be";
			when "0100110011" =>
				volume_next <= X"aa16";
			when "0100110100" =>
				volume_next <= X"aa6d";
			when "0100110101" =>
				volume_next <= X"aac5";
			when "0100110110" =>
				volume_next <= X"ab1c";
			when "0100110111" =>
				volume_next <= X"ab73";
			when "0100111000" =>
				volume_next <= X"abca";
			when "0100111001" =>
				volume_next <= X"ac20";
			when "0100111010" =>
				volume_next <= X"ac76";
			when "0100111011" =>
				volume_next <= X"accc";
			when "0100111100" =>
				volume_next <= X"ad21";
			when "0100111101" =>
				volume_next <= X"ad77";
			when "0100111110" =>
				volume_next <= X"adcb";
			when "0100111111" =>
				volume_next <= X"ae20";
			when "0101000000" =>
				volume_next <= X"ae74";
			when "0101000001" =>
				volume_next <= X"aec8";
			when "0101000010" =>
				volume_next <= X"af1c";
			when "0101000011" =>
				volume_next <= X"af70";
			when "0101000100" =>
				volume_next <= X"afc3";
			when "0101000101" =>
				volume_next <= X"b016";
			when "0101000110" =>
				volume_next <= X"b068";
			when "0101000111" =>
				volume_next <= X"b0bb";
			when "0101001000" =>
				volume_next <= X"b10d";
			when "0101001001" =>
				volume_next <= X"b15f";
			when "0101001010" =>
				volume_next <= X"b1b0";
			when "0101001011" =>
				volume_next <= X"b201";
			when "0101001100" =>
				volume_next <= X"b252";
			when "0101001101" =>
				volume_next <= X"b2a3";
			when "0101001110" =>
				volume_next <= X"b2f4";
			when "0101001111" =>
				volume_next <= X"b344";
			when "0101010000" =>
				volume_next <= X"b393";
			when "0101010001" =>
				volume_next <= X"b3e3";
			when "0101010010" =>
				volume_next <= X"b432";
			when "0101010011" =>
				volume_next <= X"b481";
			when "0101010100" =>
				volume_next <= X"b4d0";
			when "0101010101" =>
				volume_next <= X"b51f";
			when "0101010110" =>
				volume_next <= X"b56d";
			when "0101010111" =>
				volume_next <= X"b5bb";
			when "0101011000" =>
				volume_next <= X"b608";
			when "0101011001" =>
				volume_next <= X"b656";
			when "0101011010" =>
				volume_next <= X"b6a3";
			when "0101011011" =>
				volume_next <= X"b6f0";
			when "0101011100" =>
				volume_next <= X"b73c";
			when "0101011101" =>
				volume_next <= X"b789";
			when "0101011110" =>
				volume_next <= X"b7d5";
			when "0101011111" =>
				volume_next <= X"b821";
			when "0101100000" =>
				volume_next <= X"b86c";
			when "0101100001" =>
				volume_next <= X"b8b7";
			when "0101100010" =>
				volume_next <= X"b902";
			when "0101100011" =>
				volume_next <= X"b94d";
			when "0101100100" =>
				volume_next <= X"b998";
			when "0101100101" =>
				volume_next <= X"b9e2";
			when "0101100110" =>
				volume_next <= X"ba2c";
			when "0101100111" =>
				volume_next <= X"ba75";
			when "0101101000" =>
				volume_next <= X"babf";
			when "0101101001" =>
				volume_next <= X"bb08";
			when "0101101010" =>
				volume_next <= X"bb51";
			when "0101101011" =>
				volume_next <= X"bb99";
			when "0101101100" =>
				volume_next <= X"bbe2";
			when "0101101101" =>
				volume_next <= X"bc2a";
			when "0101101110" =>
				volume_next <= X"bc72";
			when "0101101111" =>
				volume_next <= X"bcb9";
			when "0101110000" =>
				volume_next <= X"bd01";
			when "0101110001" =>
				volume_next <= X"bd48";
			when "0101110010" =>
				volume_next <= X"bd8f";
			when "0101110011" =>
				volume_next <= X"bdd5";
			when "0101110100" =>
				volume_next <= X"be1b";
			when "0101110101" =>
				volume_next <= X"be62";
			when "0101110110" =>
				volume_next <= X"bea7";
			when "0101110111" =>
				volume_next <= X"beed";
			when "0101111000" =>
				volume_next <= X"bf32";
			when "0101111001" =>
				volume_next <= X"bf77";
			when "0101111010" =>
				volume_next <= X"bfbc";
			when "0101111011" =>
				volume_next <= X"c001";
			when "0101111100" =>
				volume_next <= X"c045";
			when "0101111101" =>
				volume_next <= X"c089";
			when "0101111110" =>
				volume_next <= X"c0cd";
			when "0101111111" =>
				volume_next <= X"c110";
			when "0110000000" =>
				volume_next <= X"c154";
			when "0110000001" =>
				volume_next <= X"c197";
			when "0110000010" =>
				volume_next <= X"c1d9";
			when "0110000011" =>
				volume_next <= X"c21c";
			when "0110000100" =>
				volume_next <= X"c25e";
			when "0110000101" =>
				volume_next <= X"c2a0";
			when "0110000110" =>
				volume_next <= X"c2e2";
			when "0110000111" =>
				volume_next <= X"c324";
			when "0110001000" =>
				volume_next <= X"c365";
			when "0110001001" =>
				volume_next <= X"c3a6";
			when "0110001010" =>
				volume_next <= X"c3e7";
			when "0110001011" =>
				volume_next <= X"c428";
			when "0110001100" =>
				volume_next <= X"c468";
			when "0110001101" =>
				volume_next <= X"c4a8";
			when "0110001110" =>
				volume_next <= X"c4e8";
			when "0110001111" =>
				volume_next <= X"c528";
			when "0110010000" =>
				volume_next <= X"c567";
			when "0110010001" =>
				volume_next <= X"c5a6";
			when "0110010010" =>
				volume_next <= X"c5e5";
			when "0110010011" =>
				volume_next <= X"c624";
			when "0110010100" =>
				volume_next <= X"c662";
			when "0110010101" =>
				volume_next <= X"c6a0";
			when "0110010110" =>
				volume_next <= X"c6de";
			when "0110010111" =>
				volume_next <= X"c71c";
			when "0110011000" =>
				volume_next <= X"c75a";
			when "0110011001" =>
				volume_next <= X"c797";
			when "0110011010" =>
				volume_next <= X"c7d4";
			when "0110011011" =>
				volume_next <= X"c811";
			when "0110011100" =>
				volume_next <= X"c84d";
			when "0110011101" =>
				volume_next <= X"c88a";
			when "0110011110" =>
				volume_next <= X"c8c6";
			when "0110011111" =>
				volume_next <= X"c902";
			when "0110100000" =>
				volume_next <= X"c93e";
			when "0110100001" =>
				volume_next <= X"c979";
			when "0110100010" =>
				volume_next <= X"c9b4";
			when "0110100011" =>
				volume_next <= X"c9ef";
			when "0110100100" =>
				volume_next <= X"ca2a";
			when "0110100101" =>
				volume_next <= X"ca64";
			when "0110100110" =>
				volume_next <= X"ca9f";
			when "0110100111" =>
				volume_next <= X"cad9";
			when "0110101000" =>
				volume_next <= X"cb13";
			when "0110101001" =>
				volume_next <= X"cb4c";
			when "0110101010" =>
				volume_next <= X"cb86";
			when "0110101011" =>
				volume_next <= X"cbbf";
			when "0110101100" =>
				volume_next <= X"cbf8";
			when "0110101101" =>
				volume_next <= X"cc31";
			when "0110101110" =>
				volume_next <= X"cc69";
			when "0110101111" =>
				volume_next <= X"cca1";
			when "0110110000" =>
				volume_next <= X"ccd9";
			when "0110110001" =>
				volume_next <= X"cd11";
			when "0110110010" =>
				volume_next <= X"cd49";
			when "0110110011" =>
				volume_next <= X"cd80";
			when "0110110100" =>
				volume_next <= X"cdb8";
			when "0110110101" =>
				volume_next <= X"cdee";
			when "0110110110" =>
				volume_next <= X"ce25";
			when "0110110111" =>
				volume_next <= X"ce5c";
			when "0110111000" =>
				volume_next <= X"ce92";
			when "0110111001" =>
				volume_next <= X"cec8";
			when "0110111010" =>
				volume_next <= X"cefe";
			when "0110111011" =>
				volume_next <= X"cf34";
			when "0110111100" =>
				volume_next <= X"cf69";
			when "0110111101" =>
				volume_next <= X"cf9f";
			when "0110111110" =>
				volume_next <= X"cfd4";
			when "0110111111" =>
				volume_next <= X"d008";
			when "0111000000" =>
				volume_next <= X"d03d";
			when "0111000001" =>
				volume_next <= X"d071";
			when "0111000010" =>
				volume_next <= X"d0a6";
			when "0111000011" =>
				volume_next <= X"d0da";
			when "0111000100" =>
				volume_next <= X"d10d";
			when "0111000101" =>
				volume_next <= X"d141";
			when "0111000110" =>
				volume_next <= X"d174";
			when "0111000111" =>
				volume_next <= X"d1a8";
			when "0111001000" =>
				volume_next <= X"d1db";
			when "0111001001" =>
				volume_next <= X"d20d";
			when "0111001010" =>
				volume_next <= X"d240";
			when "0111001011" =>
				volume_next <= X"d272";
			when "0111001100" =>
				volume_next <= X"d2a4";
			when "0111001101" =>
				volume_next <= X"d2d6";
			when "0111001110" =>
				volume_next <= X"d308";
			when "0111001111" =>
				volume_next <= X"d33a";
			when "0111010000" =>
				volume_next <= X"d36b";
			when "0111010001" =>
				volume_next <= X"d39c";
			when "0111010010" =>
				volume_next <= X"d3cd";
			when "0111010011" =>
				volume_next <= X"d3fe";
			when "0111010100" =>
				volume_next <= X"d42e";
			when "0111010101" =>
				volume_next <= X"d45e";
			when "0111010110" =>
				volume_next <= X"d48f";
			when "0111010111" =>
				volume_next <= X"d4bf";
			when "0111011000" =>
				volume_next <= X"d4ee";
			when "0111011001" =>
				volume_next <= X"d51e";
			when "0111011010" =>
				volume_next <= X"d54d";
			when "0111011011" =>
				volume_next <= X"d57c";
			when "0111011100" =>
				volume_next <= X"d5ab";
			when "0111011101" =>
				volume_next <= X"d5da";
			when "0111011110" =>
				volume_next <= X"d609";
			when "0111011111" =>
				volume_next <= X"d637";
			when "0111100000" =>
				volume_next <= X"d665";
			when "0111100001" =>
				volume_next <= X"d693";
			when "0111100010" =>
				volume_next <= X"d6c1";
			when "0111100011" =>
				volume_next <= X"d6ee";
			when "0111100100" =>
				volume_next <= X"d71c";
			when "0111100101" =>
				volume_next <= X"d749";
			when "0111100110" =>
				volume_next <= X"d776";
			when "0111100111" =>
				volume_next <= X"d7a3";
			when "0111101000" =>
				volume_next <= X"d7d0";
			when "0111101001" =>
				volume_next <= X"d7fc";
			when "0111101010" =>
				volume_next <= X"d828";
			when "0111101011" =>
				volume_next <= X"d854";
			when "0111101100" =>
				volume_next <= X"d880";
			when "0111101101" =>
				volume_next <= X"d8ac";
			when "0111101110" =>
				volume_next <= X"d8d8";
			when "0111101111" =>
				volume_next <= X"d903";
			when "0111110000" =>
				volume_next <= X"d92e";
			when "0111110001" =>
				volume_next <= X"d959";
			when "0111110010" =>
				volume_next <= X"d984";
			when "0111110011" =>
				volume_next <= X"d9af";
			when "0111110100" =>
				volume_next <= X"d9d9";
			when "0111110101" =>
				volume_next <= X"da03";
			when "0111110110" =>
				volume_next <= X"da2d";
			when "0111110111" =>
				volume_next <= X"da57";
			when "0111111000" =>
				volume_next <= X"da81";
			when "0111111001" =>
				volume_next <= X"daab";
			when "0111111010" =>
				volume_next <= X"dad4";
			when "0111111011" =>
				volume_next <= X"dafd";
			when "0111111100" =>
				volume_next <= X"db26";
			when "0111111101" =>
				volume_next <= X"db4f";
			when "0111111110" =>
				volume_next <= X"db78";
			when "0111111111" =>
				volume_next <= X"dba0";
			when "1000000000" =>
				volume_next <= X"dbc8";
			when "1000000001" =>
				volume_next <= X"dbf1";
			when "1000000010" =>
				volume_next <= X"dc19";
			when "1000000011" =>
				volume_next <= X"dc40";
			when "1000000100" =>
				volume_next <= X"dc68";
			when "1000000101" =>
				volume_next <= X"dc8f";
			when "1000000110" =>
				volume_next <= X"dcb7";
			when "1000000111" =>
				volume_next <= X"dcde";
			when "1000001000" =>
				volume_next <= X"dd05";
			when "1000001001" =>
				volume_next <= X"dd2c";
			when "1000001010" =>
				volume_next <= X"dd52";
			when "1000001011" =>
				volume_next <= X"dd79";
			when "1000001100" =>
				volume_next <= X"dd9f";
			when "1000001101" =>
				volume_next <= X"ddc5";
			when "1000001110" =>
				volume_next <= X"ddeb";
			when "1000001111" =>
				volume_next <= X"de11";
			when "1000010000" =>
				volume_next <= X"de36";
			when "1000010001" =>
				volume_next <= X"de5c";
			when "1000010010" =>
				volume_next <= X"de81";
			when "1000010011" =>
				volume_next <= X"dea6";
			when "1000010100" =>
				volume_next <= X"decb";
			when "1000010101" =>
				volume_next <= X"def0";
			when "1000010110" =>
				volume_next <= X"df15";
			when "1000010111" =>
				volume_next <= X"df39";
			when "1000011000" =>
				volume_next <= X"df5d";
			when "1000011001" =>
				volume_next <= X"df82";
			when "1000011010" =>
				volume_next <= X"dfa6";
			when "1000011011" =>
				volume_next <= X"dfc9";
			when "1000011100" =>
				volume_next <= X"dfed";
			when "1000011101" =>
				volume_next <= X"e011";
			when "1000011110" =>
				volume_next <= X"e034";
			when "1000011111" =>
				volume_next <= X"e057";
			when "1000100000" =>
				volume_next <= X"e07a";
			when "1000100001" =>
				volume_next <= X"e09d";
			when "1000100010" =>
				volume_next <= X"e0c0";
			when "1000100011" =>
				volume_next <= X"e0e2";
			when "1000100100" =>
				volume_next <= X"e105";
			when "1000100101" =>
				volume_next <= X"e127";
			when "1000100110" =>
				volume_next <= X"e149";
			when "1000100111" =>
				volume_next <= X"e16b";
			when "1000101000" =>
				volume_next <= X"e18d";
			when "1000101001" =>
				volume_next <= X"e1af";
			when "1000101010" =>
				volume_next <= X"e1d0";
			when "1000101011" =>
				volume_next <= X"e1f2";
			when "1000101100" =>
				volume_next <= X"e213";
			when "1000101101" =>
				volume_next <= X"e234";
			when "1000101110" =>
				volume_next <= X"e255";
			when "1000101111" =>
				volume_next <= X"e276";
			when "1000110000" =>
				volume_next <= X"e296";
			when "1000110001" =>
				volume_next <= X"e2b7";
			when "1000110010" =>
				volume_next <= X"e2d7";
			when "1000110011" =>
				volume_next <= X"e2f7";
			when "1000110100" =>
				volume_next <= X"e317";
			when "1000110101" =>
				volume_next <= X"e337";
			when "1000110110" =>
				volume_next <= X"e357";
			when "1000110111" =>
				volume_next <= X"e377";
			when "1000111000" =>
				volume_next <= X"e396";
			when "1000111001" =>
				volume_next <= X"e3b6";
			when "1000111010" =>
				volume_next <= X"e3d5";
			when "1000111011" =>
				volume_next <= X"e3f4";
			when "1000111100" =>
				volume_next <= X"e413";
			when "1000111101" =>
				volume_next <= X"e432";
			when "1000111110" =>
				volume_next <= X"e450";
			when "1000111111" =>
				volume_next <= X"e46f";
			when "1001000000" =>
				volume_next <= X"e48d";
			when "1001000001" =>
				volume_next <= X"e4ab";
			when "1001000010" =>
				volume_next <= X"e4c9";
			when "1001000011" =>
				volume_next <= X"e4e7";
			when "1001000100" =>
				volume_next <= X"e505";
			when "1001000101" =>
				volume_next <= X"e523";
			when "1001000110" =>
				volume_next <= X"e541";
			when "1001000111" =>
				volume_next <= X"e55e";
			when "1001001000" =>
				volume_next <= X"e57b";
			when "1001001001" =>
				volume_next <= X"e598";
			when "1001001010" =>
				volume_next <= X"e5b6";
			when "1001001011" =>
				volume_next <= X"e5d2";
			when "1001001100" =>
				volume_next <= X"e5ef";
			when "1001001101" =>
				volume_next <= X"e60c";
			when "1001001110" =>
				volume_next <= X"e628";
			when "1001001111" =>
				volume_next <= X"e645";
			when "1001010000" =>
				volume_next <= X"e661";
			when "1001010001" =>
				volume_next <= X"e67d";
			when "1001010010" =>
				volume_next <= X"e699";
			when "1001010011" =>
				volume_next <= X"e6b5";
			when "1001010100" =>
				volume_next <= X"e6d1";
			when "1001010101" =>
				volume_next <= X"e6ec";
			when "1001010110" =>
				volume_next <= X"e708";
			when "1001010111" =>
				volume_next <= X"e723";
			when "1001011000" =>
				volume_next <= X"e73f";
			when "1001011001" =>
				volume_next <= X"e75a";
			when "1001011010" =>
				volume_next <= X"e775";
			when "1001011011" =>
				volume_next <= X"e790";
			when "1001011100" =>
				volume_next <= X"e7aa";
			when "1001011101" =>
				volume_next <= X"e7c5";
			when "1001011110" =>
				volume_next <= X"e7e0";
			when "1001011111" =>
				volume_next <= X"e7fa";
			when "1001100000" =>
				volume_next <= X"e814";
			when "1001100001" =>
				volume_next <= X"e82f";
			when "1001100010" =>
				volume_next <= X"e849";
			when "1001100011" =>
				volume_next <= X"e862";
			when "1001100100" =>
				volume_next <= X"e87c";
			when "1001100101" =>
				volume_next <= X"e896";
			when "1001100110" =>
				volume_next <= X"e8b0";
			when "1001100111" =>
				volume_next <= X"e8c9";
			when "1001101000" =>
				volume_next <= X"e8e2";
			when "1001101001" =>
				volume_next <= X"e8fc";
			when "1001101010" =>
				volume_next <= X"e915";
			when "1001101011" =>
				volume_next <= X"e92e";
			when "1001101100" =>
				volume_next <= X"e947";
			when "1001101101" =>
				volume_next <= X"e960";
			when "1001101110" =>
				volume_next <= X"e978";
			when "1001101111" =>
				volume_next <= X"e991";
			when "1001110000" =>
				volume_next <= X"e9a9";
			when "1001110001" =>
				volume_next <= X"e9c2";
			when "1001110010" =>
				volume_next <= X"e9da";
			when "1001110011" =>
				volume_next <= X"e9f2";
			when "1001110100" =>
				volume_next <= X"ea0a";
			when "1001110101" =>
				volume_next <= X"ea22";
			when "1001110110" =>
				volume_next <= X"ea3a";
			when "1001110111" =>
				volume_next <= X"ea52";
			when "1001111000" =>
				volume_next <= X"ea69";
			when "1001111001" =>
				volume_next <= X"ea81";
			when "1001111010" =>
				volume_next <= X"ea98";
			when "1001111011" =>
				volume_next <= X"eab0";
			when "1001111100" =>
				volume_next <= X"eac7";
			when "1001111101" =>
				volume_next <= X"eade";
			when "1001111110" =>
				volume_next <= X"eaf5";
			when "1001111111" =>
				volume_next <= X"eb0c";
			when "1010000000" =>
				volume_next <= X"eb23";
			when "1010000001" =>
				volume_next <= X"eb39";
			when "1010000010" =>
				volume_next <= X"eb50";
			when "1010000011" =>
				volume_next <= X"eb66";
			when "1010000100" =>
				volume_next <= X"eb7d";
			when "1010000101" =>
				volume_next <= X"eb93";
			when "1010000110" =>
				volume_next <= X"eba9";
			when "1010000111" =>
				volume_next <= X"ebbf";
			when "1010001000" =>
				volume_next <= X"ebd6";
			when "1010001001" =>
				volume_next <= X"ebeb";
			when "1010001010" =>
				volume_next <= X"ec01";
			when "1010001011" =>
				volume_next <= X"ec17";
			when "1010001100" =>
				volume_next <= X"ec2d";
			when "1010001101" =>
				volume_next <= X"ec42";
			when "1010001110" =>
				volume_next <= X"ec58";
			when "1010001111" =>
				volume_next <= X"ec6d";
			when "1010010000" =>
				volume_next <= X"ec82";
			when "1010010001" =>
				volume_next <= X"ec98";
			when "1010010010" =>
				volume_next <= X"ecad";
			when "1010010011" =>
				volume_next <= X"ecc2";
			when "1010010100" =>
				volume_next <= X"ecd7";
			when "1010010101" =>
				volume_next <= X"eceb";
			when "1010010110" =>
				volume_next <= X"ed00";
			when "1010010111" =>
				volume_next <= X"ed15";
			when "1010011000" =>
				volume_next <= X"ed29";
			when "1010011001" =>
				volume_next <= X"ed3e";
			when "1010011010" =>
				volume_next <= X"ed52";
			when "1010011011" =>
				volume_next <= X"ed67";
			when "1010011100" =>
				volume_next <= X"ed7b";
			when "1010011101" =>
				volume_next <= X"ed8f";
			when "1010011110" =>
				volume_next <= X"eda3";
			when "1010011111" =>
				volume_next <= X"edb7";
			when "1010100000" =>
				volume_next <= X"edcb";
			when "1010100001" =>
				volume_next <= X"eddf";
			when "1010100010" =>
				volume_next <= X"edf3";
			when "1010100011" =>
				volume_next <= X"ee06";
			when "1010100100" =>
				volume_next <= X"ee1a";
			when "1010100101" =>
				volume_next <= X"ee2d";
			when "1010100110" =>
				volume_next <= X"ee41";
			when "1010100111" =>
				volume_next <= X"ee54";
			when "1010101000" =>
				volume_next <= X"ee67";
			when "1010101001" =>
				volume_next <= X"ee7b";
			when "1010101010" =>
				volume_next <= X"ee8e";
			when "1010101011" =>
				volume_next <= X"eea1";
			when "1010101100" =>
				volume_next <= X"eeb4";
			when "1010101101" =>
				volume_next <= X"eec7";
			when "1010101110" =>
				volume_next <= X"eed9";
			when "1010101111" =>
				volume_next <= X"eeec";
			when "1010110000" =>
				volume_next <= X"eeff";
			when "1010110001" =>
				volume_next <= X"ef11";
			when "1010110010" =>
				volume_next <= X"ef24";
			when "1010110011" =>
				volume_next <= X"ef36";
			when "1010110100" =>
				volume_next <= X"ef49";
			when "1010110101" =>
				volume_next <= X"ef5b";
			when "1010110110" =>
				volume_next <= X"ef6d";
			when "1010110111" =>
				volume_next <= X"ef80";
			when "1010111000" =>
				volume_next <= X"ef92";
			when "1010111001" =>
				volume_next <= X"efa4";
			when "1010111010" =>
				volume_next <= X"efb6";
			when "1010111011" =>
				volume_next <= X"efc8";
			when "1010111100" =>
				volume_next <= X"efda";
			when "1010111101" =>
				volume_next <= X"efeb";
			when "1010111110" =>
				volume_next <= X"effd";
			when "1010111111" =>
				volume_next <= X"f00f";
			when "1011000000" =>
				volume_next <= X"f020";
			when "1011000001" =>
				volume_next <= X"f032";
			when "1011000010" =>
				volume_next <= X"f043";
			when "1011000011" =>
				volume_next <= X"f055";
			when "1011000100" =>
				volume_next <= X"f066";
			when "1011000101" =>
				volume_next <= X"f077";
			when "1011000110" =>
				volume_next <= X"f089";
			when "1011000111" =>
				volume_next <= X"f09a";
			when "1011001000" =>
				volume_next <= X"f0ab";
			when "1011001001" =>
				volume_next <= X"f0bc";
			when "1011001010" =>
				volume_next <= X"f0cd";
			when "1011001011" =>
				volume_next <= X"f0de";
			when "1011001100" =>
				volume_next <= X"f0ef";
			when "1011001101" =>
				volume_next <= X"f100";
			when "1011001110" =>
				volume_next <= X"f110";
			when "1011001111" =>
				volume_next <= X"f121";
			when "1011010000" =>
				volume_next <= X"f132";
			when "1011010001" =>
				volume_next <= X"f142";
			when "1011010010" =>
				volume_next <= X"f153";
			when "1011010011" =>
				volume_next <= X"f163";
			when "1011010100" =>
				volume_next <= X"f174";
			when "1011010101" =>
				volume_next <= X"f184";
			when "1011010110" =>
				volume_next <= X"f195";
			when "1011010111" =>
				volume_next <= X"f1a5";
			when "1011011000" =>
				volume_next <= X"f1b5";
			when "1011011001" =>
				volume_next <= X"f1c5";
			when "1011011010" =>
				volume_next <= X"f1d6";
			when "1011011011" =>
				volume_next <= X"f1e6";
			when "1011011100" =>
				volume_next <= X"f1f6";
			when "1011011101" =>
				volume_next <= X"f206";
			when "1011011110" =>
				volume_next <= X"f216";
			when "1011011111" =>
				volume_next <= X"f226";
			when "1011100000" =>
				volume_next <= X"f236";
			when "1011100001" =>
				volume_next <= X"f245";
			when "1011100010" =>
				volume_next <= X"f255";
			when "1011100011" =>
				volume_next <= X"f265";
			when "1011100100" =>
				volume_next <= X"f275";
			when "1011100101" =>
				volume_next <= X"f284";
			when "1011100110" =>
				volume_next <= X"f294";
			when "1011100111" =>
				volume_next <= X"f2a4";
			when "1011101000" =>
				volume_next <= X"f2b3";
			when "1011101001" =>
				volume_next <= X"f2c3";
			when "1011101010" =>
				volume_next <= X"f2d2";
			when "1011101011" =>
				volume_next <= X"f2e1";
			when "1011101100" =>
				volume_next <= X"f2f1";
			when "1011101101" =>
				volume_next <= X"f300";
			when "1011101110" =>
				volume_next <= X"f310";
			when "1011101111" =>
				volume_next <= X"f31f";
			when "1011110000" =>
				volume_next <= X"f32e";
			when "1011110001" =>
				volume_next <= X"f33d";
			when "1011110010" =>
				volume_next <= X"f34c";
			when "1011110011" =>
				volume_next <= X"f35c";
			when "1011110100" =>
				volume_next <= X"f36b";
			when "1011110101" =>
				volume_next <= X"f37a";
			when "1011110110" =>
				volume_next <= X"f389";
			when "1011110111" =>
				volume_next <= X"f398";
			when "1011111000" =>
				volume_next <= X"f3a7";
			when "1011111001" =>
				volume_next <= X"f3b6";
			when "1011111010" =>
				volume_next <= X"f3c5";
			when "1011111011" =>
				volume_next <= X"f3d4";
			when "1011111100" =>
				volume_next <= X"f3e2";
			when "1011111101" =>
				volume_next <= X"f3f1";
			when "1011111110" =>
				volume_next <= X"f400";
			when "1011111111" =>
				volume_next <= X"f40f";
			when "1100000000" =>
				volume_next <= X"f41e";
			when "1100000001" =>
				volume_next <= X"f42c";
			when "1100000010" =>
				volume_next <= X"f43b";
			when "1100000011" =>
				volume_next <= X"f44a";
			when "1100000100" =>
				volume_next <= X"f458";
			when "1100000101" =>
				volume_next <= X"f467";
			when "1100000110" =>
				volume_next <= X"f476";
			when "1100000111" =>
				volume_next <= X"f484";
			when "1100001000" =>
				volume_next <= X"f493";
			when "1100001001" =>
				volume_next <= X"f4a1";
			when "1100001010" =>
				volume_next <= X"f4b0";
			when "1100001011" =>
				volume_next <= X"f4be";
			when "1100001100" =>
				volume_next <= X"f4cd";
			when "1100001101" =>
				volume_next <= X"f4db";
			when "1100001110" =>
				volume_next <= X"f4ea";
			when "1100001111" =>
				volume_next <= X"f4f8";
			when "1100010000" =>
				volume_next <= X"f507";
			when "1100010001" =>
				volume_next <= X"f515";
			when "1100010010" =>
				volume_next <= X"f524";
			when "1100010011" =>
				volume_next <= X"f532";
			when "1100010100" =>
				volume_next <= X"f540";
			when "1100010101" =>
				volume_next <= X"f54f";
			when "1100010110" =>
				volume_next <= X"f55d";
			when "1100010111" =>
				volume_next <= X"f56b";
			when "1100011000" =>
				volume_next <= X"f57a";
			when "1100011001" =>
				volume_next <= X"f588";
			when "1100011010" =>
				volume_next <= X"f596";
			when "1100011011" =>
				volume_next <= X"f5a4";
			when "1100011100" =>
				volume_next <= X"f5b3";
			when "1100011101" =>
				volume_next <= X"f5c1";
			when "1100011110" =>
				volume_next <= X"f5cf";
			when "1100011111" =>
				volume_next <= X"f5dd";
			when "1100100000" =>
				volume_next <= X"f5ec";
			when "1100100001" =>
				volume_next <= X"f5fa";
			when "1100100010" =>
				volume_next <= X"f608";
			when "1100100011" =>
				volume_next <= X"f616";
			when "1100100100" =>
				volume_next <= X"f624";
			when "1100100101" =>
				volume_next <= X"f633";
			when "1100100110" =>
				volume_next <= X"f641";
			when "1100100111" =>
				volume_next <= X"f64f";
			when "1100101000" =>
				volume_next <= X"f65d";
			when "1100101001" =>
				volume_next <= X"f66b";
			when "1100101010" =>
				volume_next <= X"f67a";
			when "1100101011" =>
				volume_next <= X"f688";
			when "1100101100" =>
				volume_next <= X"f696";
			when "1100101101" =>
				volume_next <= X"f6a4";
			when "1100101110" =>
				volume_next <= X"f6b2";
			when "1100101111" =>
				volume_next <= X"f6c0";
			when "1100110000" =>
				volume_next <= X"f6cf";
			when "1100110001" =>
				volume_next <= X"f6dd";
			when "1100110010" =>
				volume_next <= X"f6eb";
			when "1100110011" =>
				volume_next <= X"f6f9";
			when "1100110100" =>
				volume_next <= X"f707";
			when "1100110101" =>
				volume_next <= X"f716";
			when "1100110110" =>
				volume_next <= X"f724";
			when "1100110111" =>
				volume_next <= X"f732";
			when "1100111000" =>
				volume_next <= X"f740";
			when "1100111001" =>
				volume_next <= X"f74e";
			when "1100111010" =>
				volume_next <= X"f75d";
			when "1100111011" =>
				volume_next <= X"f76b";
			when "1100111100" =>
				volume_next <= X"f779";
			when "1100111101" =>
				volume_next <= X"f787";
			when "1100111110" =>
				volume_next <= X"f796";
			when "1100111111" =>
				volume_next <= X"f7a4";
			when "1101000000" =>
				volume_next <= X"f7b2";
			when "1101000001" =>
				volume_next <= X"f7c0";
			when "1101000010" =>
				volume_next <= X"f7cf";
			when "1101000011" =>
				volume_next <= X"f7dd";
			when "1101000100" =>
				volume_next <= X"f7eb";
			when "1101000101" =>
				volume_next <= X"f7fa";
			when "1101000110" =>
				volume_next <= X"f808";
			when "1101000111" =>
				volume_next <= X"f817";
			when "1101001000" =>
				volume_next <= X"f825";
			when "1101001001" =>
				volume_next <= X"f833";
			when "1101001010" =>
				volume_next <= X"f842";
			when "1101001011" =>
				volume_next <= X"f850";
			when "1101001100" =>
				volume_next <= X"f85f";
			when "1101001101" =>
				volume_next <= X"f86d";
			when "1101001110" =>
				volume_next <= X"f87c";
			when "1101001111" =>
				volume_next <= X"f88a";
			when "1101010000" =>
				volume_next <= X"f899";
			when "1101010001" =>
				volume_next <= X"f8a7";
			when "1101010010" =>
				volume_next <= X"f8b6";
			when "1101010011" =>
				volume_next <= X"f8c4";
			when "1101010100" =>
				volume_next <= X"f8d3";
			when "1101010101" =>
				volume_next <= X"f8e2";
			when "1101010110" =>
				volume_next <= X"f8f0";
			when "1101010111" =>
				volume_next <= X"f8ff";
			when "1101011000" =>
				volume_next <= X"f90e";
			when "1101011001" =>
				volume_next <= X"f91d";
			when "1101011010" =>
				volume_next <= X"f92b";
			when "1101011011" =>
				volume_next <= X"f93a";
			when "1101011100" =>
				volume_next <= X"f949";
			when "1101011101" =>
				volume_next <= X"f958";
			when "1101011110" =>
				volume_next <= X"f967";
			when "1101011111" =>
				volume_next <= X"f976";
			when "1101100000" =>
				volume_next <= X"f984";
			when "1101100001" =>
				volume_next <= X"f993";
			when "1101100010" =>
				volume_next <= X"f9a2";
			when "1101100011" =>
				volume_next <= X"f9b1";
			when "1101100100" =>
				volume_next <= X"f9c1";
			when "1101100101" =>
				volume_next <= X"f9d0";
			when "1101100110" =>
				volume_next <= X"f9df";
			when "1101100111" =>
				volume_next <= X"f9ee";
			when "1101101000" =>
				volume_next <= X"f9fd";
			when "1101101001" =>
				volume_next <= X"fa0c";
			when "1101101010" =>
				volume_next <= X"fa1c";
			when "1101101011" =>
				volume_next <= X"fa2b";
			when "1101101100" =>
				volume_next <= X"fa3a";
			when "1101101101" =>
				volume_next <= X"fa4a";
			when "1101101110" =>
				volume_next <= X"fa59";
			when "1101101111" =>
				volume_next <= X"fa68";
			when "1101110000" =>
				volume_next <= X"fa78";
			when "1101110001" =>
				volume_next <= X"fa87";
			when "1101110010" =>
				volume_next <= X"fa97";
			when "1101110011" =>
				volume_next <= X"faa7";
			when "1101110100" =>
				volume_next <= X"fab6";
			when "1101110101" =>
				volume_next <= X"fac6";
			when "1101110110" =>
				volume_next <= X"fad6";
			when "1101110111" =>
				volume_next <= X"fae5";
			when "1101111000" =>
				volume_next <= X"faf5";
			when "1101111001" =>
				volume_next <= X"fb05";
			when "1101111010" =>
				volume_next <= X"fb15";
			when "1101111011" =>
				volume_next <= X"fb25";
			when "1101111100" =>
				volume_next <= X"fb35";
			when "1101111101" =>
				volume_next <= X"fb45";
			when "1101111110" =>
				volume_next <= X"fb55";
			when "1101111111" =>
				volume_next <= X"fb65";
			when "1110000000" =>
				volume_next <= X"fb75";
			when "1110000001" =>
				volume_next <= X"fb86";
			when "1110000010" =>
				volume_next <= X"fb96";
			when "1110000011" =>
				volume_next <= X"fba6";
			when "1110000100" =>
				volume_next <= X"fbb7";
			when "1110000101" =>
				volume_next <= X"fbc7";
			when "1110000110" =>
				volume_next <= X"fbd7";
			when "1110000111" =>
				volume_next <= X"fbe8";
			when "1110001000" =>
				volume_next <= X"fbf9";
			when "1110001001" =>
				volume_next <= X"fc09";
			when "1110001010" =>
				volume_next <= X"fc1a";
			when "1110001011" =>
				volume_next <= X"fc2b";
			when "1110001100" =>
				volume_next <= X"fc3b";
			when "1110001101" =>
				volume_next <= X"fc4c";
			when "1110001110" =>
				volume_next <= X"fc5d";
			when "1110001111" =>
				volume_next <= X"fc6e";
			when "1110010000" =>
				volume_next <= X"fc7f";
			when "1110010001" =>
				volume_next <= X"fc90";
			when "1110010010" =>
				volume_next <= X"fca1";
			when "1110010011" =>
				volume_next <= X"fcb3";
			when "1110010100" =>
				volume_next <= X"fcc4";
			when "1110010101" =>
				volume_next <= X"fcd5";
			when "1110010110" =>
				volume_next <= X"fce6";
			when "1110010111" =>
				volume_next <= X"fcf8";
			when "1110011000" =>
				volume_next <= X"fd09";
			when "1110011001" =>
				volume_next <= X"fd1b";
			when "1110011010" =>
				volume_next <= X"fd2d";
			when "1110011011" =>
				volume_next <= X"fd3e";
			when "1110011100" =>
				volume_next <= X"fd50";
			when "1110011101" =>
				volume_next <= X"fd62";
			when "1110011110" =>
				volume_next <= X"fd74";
			when "1110011111" =>
				volume_next <= X"fd86";
			when "1110100000" =>
				volume_next <= X"fd98";
			when "1110100001" =>
				volume_next <= X"fdaa";
			when "1110100010" =>
				volume_next <= X"fdbc";
			when "1110100011" =>
				volume_next <= X"fdce";
			when "1110100100" =>
				volume_next <= X"fde0";
			when "1110100101" =>
				volume_next <= X"fdf3";
			when "1110100110" =>
				volume_next <= X"fe05";
			when "1110100111" =>
				volume_next <= X"fe18";
			when "1110101000" =>
				volume_next <= X"fe2a";
			when "1110101001" =>
				volume_next <= X"fe3d";
			when "1110101010" =>
				volume_next <= X"fe50";
			when "1110101011" =>
				volume_next <= X"fe62";
			when "1110101100" =>
				volume_next <= X"fe75";
			when "1110101101" =>
				volume_next <= X"fe88";
			when "1110101110" =>
				volume_next <= X"fe9b";
			when "1110101111" =>
				volume_next <= X"feae";
			when "1110110000" =>
				volume_next <= X"fec1";
			when "1110110001" =>
				volume_next <= X"fed5";
			when "1110110010" =>
				volume_next <= X"fee8";
			when "1110110011" =>
				volume_next <= X"fefb";
			when "1110110100" =>
				volume_next <= X"ff0f";
			when "1110110101" =>
				volume_next <= X"ff22";
			when "1110110110" =>
				volume_next <= X"ff36";
			when "1110110111" =>
				volume_next <= X"ff4a";
			when "1110111000" =>
				volume_next <= X"ff5d";
			when "1110111001" =>
				volume_next <= X"ff71";
			when "1110111010" =>
				volume_next <= X"ff85";
			when "1110111011" =>
				volume_next <= X"ff99";
			when "1110111100" =>
				volume_next <= X"ffad";
			when "1110111101" =>
				volume_next <= X"ffc1";
			when "1110111110" =>
				volume_next <= X"ffd6";
			when "1110111111" =>
				volume_next <= X"ffea";
			when "1111000000" =>
				volume_next <= X"ffff";
			when others =>
				volume_next <= X"ffff";
		end case;
        end process;

	-- output
	volume_out <= volume_reg;
		
END vhdl;
